// Copyright Copyright Fraunhofer Institute for Applied and Integrated Security (AISEC).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

$fwrite(f,"----------------------------------------------------------------\n");   
$fwrite(f,"-- PQ Pointwise-Multiplication (Falcon-1024)\n");
$fwrite(f,"----------------------------------------------------------------\n");   
     
// Write IMEM from File
write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq_mul_falcon-1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- IMEM\n");
// Read IMEM  
for (int i=0 ; i<129 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end     

 // Write DMEM from File
write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq_mul_falcon-1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- DMEM\n");
// Read DMEM  
for (int i=0 ; i<16 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end   
	   
$fwrite(f,"----------------------------------------------------------------\n");   

// Set Instruction Counter to zero (optional)
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );

// Start Programm in IMEM
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(CmdExecute), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
cc_start = cc;
// Poll on Status Register until Programm is finished
rdbk = '1;
while (rdbk != '0) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
end 

// Measure CC
cc_stop = cc; 
cc_count_falcon1024_pointwise_mul = cc_stop - cc_start;        
       
// Read DMEM  
for (int i=0 ; i<1024 ; i++) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+128), .tl_o(tl_o), .tl_i(tl_i_d) );
    
    case(i)
	0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	5   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	6   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	7   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	8   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	9   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	10   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	11   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	12   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	13   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	14   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	15   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	16   :   assert (rdbk == 32'd256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	17   :   assert (rdbk == 32'd289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	18   :   assert (rdbk == 32'd324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	19   :   assert (rdbk == 32'd361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	20   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	21   :   assert (rdbk == 32'd441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	22   :   assert (rdbk == 32'd484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	23   :   assert (rdbk == 32'd529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	24   :   assert (rdbk == 32'd576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	25   :   assert (rdbk == 32'd625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	26   :   assert (rdbk == 32'd676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	27   :   assert (rdbk == 32'd729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	28   :   assert (rdbk == 32'd784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	29   :   assert (rdbk == 32'd841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	30   :   assert (rdbk == 32'd900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	31   :   assert (rdbk == 32'd961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	32   :   assert (rdbk == 32'd1024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	33   :   assert (rdbk == 32'd1089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	34   :   assert (rdbk == 32'd1156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	35   :   assert (rdbk == 32'd1225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	36   :   assert (rdbk == 32'd1296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	37   :   assert (rdbk == 32'd1369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	38   :   assert (rdbk == 32'd1444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	39   :   assert (rdbk == 32'd1521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	40   :   assert (rdbk == 32'd1600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	41   :   assert (rdbk == 32'd1681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	42   :   assert (rdbk == 32'd1764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	43   :   assert (rdbk == 32'd1849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	44   :   assert (rdbk == 32'd1936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	45   :   assert (rdbk == 32'd2025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	46   :   assert (rdbk == 32'd2116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	47   :   assert (rdbk == 32'd2209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	48   :   assert (rdbk == 32'd2304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	49   :   assert (rdbk == 32'd2401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	50   :   assert (rdbk == 32'd2500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	51   :   assert (rdbk == 32'd2601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	52   :   assert (rdbk == 32'd2704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	53   :   assert (rdbk == 32'd2809) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	54   :   assert (rdbk == 32'd2916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	55   :   assert (rdbk == 32'd3025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	56   :   assert (rdbk == 32'd3136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	57   :   assert (rdbk == 32'd3249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	58   :   assert (rdbk == 32'd3364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	59   :   assert (rdbk == 32'd3481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	60   :   assert (rdbk == 32'd3600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	61   :   assert (rdbk == 32'd3721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	62   :   assert (rdbk == 32'd3844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	63   :   assert (rdbk == 32'd3969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	64   :   assert (rdbk == 32'd4096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	65   :   assert (rdbk == 32'd4225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	66   :   assert (rdbk == 32'd4356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	67   :   assert (rdbk == 32'd4489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	68   :   assert (rdbk == 32'd4624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	69   :   assert (rdbk == 32'd4761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	70   :   assert (rdbk == 32'd4900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	71   :   assert (rdbk == 32'd5041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	72   :   assert (rdbk == 32'd5184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	73   :   assert (rdbk == 32'd5329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	74   :   assert (rdbk == 32'd5476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	75   :   assert (rdbk == 32'd5625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	76   :   assert (rdbk == 32'd5776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	77   :   assert (rdbk == 32'd5929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	78   :   assert (rdbk == 32'd6084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	79   :   assert (rdbk == 32'd6241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	80   :   assert (rdbk == 32'd6400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	81   :   assert (rdbk == 32'd6561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	82   :   assert (rdbk == 32'd6724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	83   :   assert (rdbk == 32'd6889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	84   :   assert (rdbk == 32'd7056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	85   :   assert (rdbk == 32'd7225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	86   :   assert (rdbk == 32'd7396) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	87   :   assert (rdbk == 32'd7569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	88   :   assert (rdbk == 32'd7744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	89   :   assert (rdbk == 32'd7921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	90   :   assert (rdbk == 32'd8100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	91   :   assert (rdbk == 32'd8281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	92   :   assert (rdbk == 32'd8464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	93   :   assert (rdbk == 32'd8649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	94   :   assert (rdbk == 32'd8836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	95   :   assert (rdbk == 32'd9025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	96   :   assert (rdbk == 32'd9216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	97   :   assert (rdbk == 32'd9409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	98   :   assert (rdbk == 32'd9604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	99   :   assert (rdbk == 32'd9801) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	100   :   assert (rdbk == 32'd10000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	101   :   assert (rdbk == 32'd10201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	102   :   assert (rdbk == 32'd10404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	103   :   assert (rdbk == 32'd10609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	104   :   assert (rdbk == 32'd10816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	105   :   assert (rdbk == 32'd11025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	106   :   assert (rdbk == 32'd11236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	107   :   assert (rdbk == 32'd11449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	108   :   assert (rdbk == 32'd11664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	109   :   assert (rdbk == 32'd11881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	110   :   assert (rdbk == 32'd12100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	111   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	112   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	113   :   assert (rdbk == 32'd480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	114   :   assert (rdbk == 32'd707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	115   :   assert (rdbk == 32'd936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	116   :   assert (rdbk == 32'd1167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	117   :   assert (rdbk == 32'd1400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	118   :   assert (rdbk == 32'd1635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	119   :   assert (rdbk == 32'd1872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	120   :   assert (rdbk == 32'd2111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	121   :   assert (rdbk == 32'd2352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	122   :   assert (rdbk == 32'd2595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	123   :   assert (rdbk == 32'd2840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	124   :   assert (rdbk == 32'd3087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	125   :   assert (rdbk == 32'd3336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	126   :   assert (rdbk == 32'd3587) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	127   :   assert (rdbk == 32'd3840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	128   :   assert (rdbk == 32'd4095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	129   :   assert (rdbk == 32'd4352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	130   :   assert (rdbk == 32'd4611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	131   :   assert (rdbk == 32'd4872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	132   :   assert (rdbk == 32'd5135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	133   :   assert (rdbk == 32'd5400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	134   :   assert (rdbk == 32'd5667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	135   :   assert (rdbk == 32'd5936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	136   :   assert (rdbk == 32'd6207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	137   :   assert (rdbk == 32'd6480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	138   :   assert (rdbk == 32'd6755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	139   :   assert (rdbk == 32'd7032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	140   :   assert (rdbk == 32'd7311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	141   :   assert (rdbk == 32'd7592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	142   :   assert (rdbk == 32'd7875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	143   :   assert (rdbk == 32'd8160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	144   :   assert (rdbk == 32'd8447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	145   :   assert (rdbk == 32'd8736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	146   :   assert (rdbk == 32'd9027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	147   :   assert (rdbk == 32'd9320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	148   :   assert (rdbk == 32'd9615) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	149   :   assert (rdbk == 32'd9912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	150   :   assert (rdbk == 32'd10211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	151   :   assert (rdbk == 32'd10512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	152   :   assert (rdbk == 32'd10815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	153   :   assert (rdbk == 32'd11120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	154   :   assert (rdbk == 32'd11427) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	155   :   assert (rdbk == 32'd11736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	156   :   assert (rdbk == 32'd12047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	157   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	158   :   assert (rdbk == 32'd386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	159   :   assert (rdbk == 32'd703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	160   :   assert (rdbk == 32'd1022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	161   :   assert (rdbk == 32'd1343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	162   :   assert (rdbk == 32'd1666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	163   :   assert (rdbk == 32'd1991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	164   :   assert (rdbk == 32'd2318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	165   :   assert (rdbk == 32'd2647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	166   :   assert (rdbk == 32'd2978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	167   :   assert (rdbk == 32'd3311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	168   :   assert (rdbk == 32'd3646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	169   :   assert (rdbk == 32'd3983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	170   :   assert (rdbk == 32'd4322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	171   :   assert (rdbk == 32'd4663) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	172   :   assert (rdbk == 32'd5006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	173   :   assert (rdbk == 32'd5351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	174   :   assert (rdbk == 32'd5698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	175   :   assert (rdbk == 32'd6047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	176   :   assert (rdbk == 32'd6398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	177   :   assert (rdbk == 32'd6751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	178   :   assert (rdbk == 32'd7106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	179   :   assert (rdbk == 32'd7463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	180   :   assert (rdbk == 32'd7822) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	181   :   assert (rdbk == 32'd8183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	182   :   assert (rdbk == 32'd8546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	183   :   assert (rdbk == 32'd8911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	184   :   assert (rdbk == 32'd9278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	185   :   assert (rdbk == 32'd9647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	186   :   assert (rdbk == 32'd10018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	187   :   assert (rdbk == 32'd10391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	188   :   assert (rdbk == 32'd10766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	189   :   assert (rdbk == 32'd11143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	190   :   assert (rdbk == 32'd11522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	191   :   assert (rdbk == 32'd11903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	192   :   assert (rdbk == 32'd12286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	193   :   assert (rdbk == 32'd382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	194   :   assert (rdbk == 32'd769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	195   :   assert (rdbk == 32'd1158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	196   :   assert (rdbk == 32'd1549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	197   :   assert (rdbk == 32'd1942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	198   :   assert (rdbk == 32'd2337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	199   :   assert (rdbk == 32'd2734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	200   :   assert (rdbk == 32'd3133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	201   :   assert (rdbk == 32'd3534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	202   :   assert (rdbk == 32'd3937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	203   :   assert (rdbk == 32'd4342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	204   :   assert (rdbk == 32'd4749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	205   :   assert (rdbk == 32'd5158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	206   :   assert (rdbk == 32'd5569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	207   :   assert (rdbk == 32'd5982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	208   :   assert (rdbk == 32'd6397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	209   :   assert (rdbk == 32'd6814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	210   :   assert (rdbk == 32'd7233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	211   :   assert (rdbk == 32'd7654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	212   :   assert (rdbk == 32'd8077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	213   :   assert (rdbk == 32'd8502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	214   :   assert (rdbk == 32'd8929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	215   :   assert (rdbk == 32'd9358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	216   :   assert (rdbk == 32'd9789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	217   :   assert (rdbk == 32'd10222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	218   :   assert (rdbk == 32'd10657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	219   :   assert (rdbk == 32'd11094) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	220   :   assert (rdbk == 32'd11533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	221   :   assert (rdbk == 32'd11974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	222   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	223   :   assert (rdbk == 32'd573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	224   :   assert (rdbk == 32'd1020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	225   :   assert (rdbk == 32'd1469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	226   :   assert (rdbk == 32'd1920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	227   :   assert (rdbk == 32'd2373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	228   :   assert (rdbk == 32'd2828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	229   :   assert (rdbk == 32'd3285) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	230   :   assert (rdbk == 32'd3744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	231   :   assert (rdbk == 32'd4205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	232   :   assert (rdbk == 32'd4668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	233   :   assert (rdbk == 32'd5133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	234   :   assert (rdbk == 32'd5600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	235   :   assert (rdbk == 32'd6069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	236   :   assert (rdbk == 32'd6540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	237   :   assert (rdbk == 32'd7013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	238   :   assert (rdbk == 32'd7488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	239   :   assert (rdbk == 32'd7965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	240   :   assert (rdbk == 32'd8444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	241   :   assert (rdbk == 32'd8925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	242   :   assert (rdbk == 32'd9408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	243   :   assert (rdbk == 32'd9893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	244   :   assert (rdbk == 32'd10380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	245   :   assert (rdbk == 32'd10869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	246   :   assert (rdbk == 32'd11360) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	247   :   assert (rdbk == 32'd11853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	248   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	249   :   assert (rdbk == 32'd556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	250   :   assert (rdbk == 32'd1055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	251   :   assert (rdbk == 32'd1556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	252   :   assert (rdbk == 32'd2059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	253   :   assert (rdbk == 32'd2564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	254   :   assert (rdbk == 32'd3071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	255   :   assert (rdbk == 32'd3580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	256   :   assert (rdbk == 32'd4091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	257   :   assert (rdbk == 32'd4604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	258   :   assert (rdbk == 32'd5119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	259   :   assert (rdbk == 32'd5636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	260   :   assert (rdbk == 32'd6155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	261   :   assert (rdbk == 32'd6676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	262   :   assert (rdbk == 32'd7199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	263   :   assert (rdbk == 32'd7724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	264   :   assert (rdbk == 32'd8251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	265   :   assert (rdbk == 32'd8780) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	266   :   assert (rdbk == 32'd9311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	267   :   assert (rdbk == 32'd9844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	268   :   assert (rdbk == 32'd10379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	269   :   assert (rdbk == 32'd10916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	270   :   assert (rdbk == 32'd11455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	271   :   assert (rdbk == 32'd11996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	272   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	273   :   assert (rdbk == 32'd795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	274   :   assert (rdbk == 32'd1342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	275   :   assert (rdbk == 32'd1891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	276   :   assert (rdbk == 32'd2442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	277   :   assert (rdbk == 32'd2995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	278   :   assert (rdbk == 32'd3550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	279   :   assert (rdbk == 32'd4107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	280   :   assert (rdbk == 32'd4666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	281   :   assert (rdbk == 32'd5227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	282   :   assert (rdbk == 32'd5790) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	283   :   assert (rdbk == 32'd6355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	284   :   assert (rdbk == 32'd6922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	285   :   assert (rdbk == 32'd7491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	286   :   assert (rdbk == 32'd8062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	287   :   assert (rdbk == 32'd8635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	288   :   assert (rdbk == 32'd9210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	289   :   assert (rdbk == 32'd9787) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	290   :   assert (rdbk == 32'd10366) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	291   :   assert (rdbk == 32'd10947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	292   :   assert (rdbk == 32'd11530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	293   :   assert (rdbk == 32'd12115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	294   :   assert (rdbk == 32'd413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	295   :   assert (rdbk == 32'd1002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	296   :   assert (rdbk == 32'd1593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	297   :   assert (rdbk == 32'd2186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	298   :   assert (rdbk == 32'd2781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	299   :   assert (rdbk == 32'd3378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	300   :   assert (rdbk == 32'd3977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	301   :   assert (rdbk == 32'd4578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	302   :   assert (rdbk == 32'd5181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	303   :   assert (rdbk == 32'd5786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	304   :   assert (rdbk == 32'd6393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	305   :   assert (rdbk == 32'd7002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	306   :   assert (rdbk == 32'd7613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	307   :   assert (rdbk == 32'd8226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	308   :   assert (rdbk == 32'd8841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	309   :   assert (rdbk == 32'd9458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	310   :   assert (rdbk == 32'd10077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	311   :   assert (rdbk == 32'd10698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	312   :   assert (rdbk == 32'd11321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	313   :   assert (rdbk == 32'd11946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	314   :   assert (rdbk == 32'd284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	315   :   assert (rdbk == 32'd913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	316   :   assert (rdbk == 32'd1544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	317   :   assert (rdbk == 32'd2177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	318   :   assert (rdbk == 32'd2812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	319   :   assert (rdbk == 32'd3449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	320   :   assert (rdbk == 32'd4088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	321   :   assert (rdbk == 32'd4729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	322   :   assert (rdbk == 32'd5372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	323   :   assert (rdbk == 32'd6017) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	324   :   assert (rdbk == 32'd6664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	325   :   assert (rdbk == 32'd7313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	326   :   assert (rdbk == 32'd7964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	327   :   assert (rdbk == 32'd8617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	328   :   assert (rdbk == 32'd9272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	329   :   assert (rdbk == 32'd9929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	330   :   assert (rdbk == 32'd10588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	331   :   assert (rdbk == 32'd11249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	332   :   assert (rdbk == 32'd11912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	333   :   assert (rdbk == 32'd288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	334   :   assert (rdbk == 32'd955) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	335   :   assert (rdbk == 32'd1624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	336   :   assert (rdbk == 32'd2295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	337   :   assert (rdbk == 32'd2968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	338   :   assert (rdbk == 32'd3643) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	339   :   assert (rdbk == 32'd4320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	340   :   assert (rdbk == 32'd4999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	341   :   assert (rdbk == 32'd5680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	342   :   assert (rdbk == 32'd6363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	343   :   assert (rdbk == 32'd7048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	344   :   assert (rdbk == 32'd7735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	345   :   assert (rdbk == 32'd8424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	346   :   assert (rdbk == 32'd9115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	347   :   assert (rdbk == 32'd9808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	348   :   assert (rdbk == 32'd10503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	349   :   assert (rdbk == 32'd11200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	350   :   assert (rdbk == 32'd11899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	351   :   assert (rdbk == 32'd311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	352   :   assert (rdbk == 32'd1014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	353   :   assert (rdbk == 32'd1719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	354   :   assert (rdbk == 32'd2426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	355   :   assert (rdbk == 32'd3135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	356   :   assert (rdbk == 32'd3846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	357   :   assert (rdbk == 32'd4559) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	358   :   assert (rdbk == 32'd5274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	359   :   assert (rdbk == 32'd5991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	360   :   assert (rdbk == 32'd6710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	361   :   assert (rdbk == 32'd7431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	362   :   assert (rdbk == 32'd8154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	363   :   assert (rdbk == 32'd8879) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	364   :   assert (rdbk == 32'd9606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	365   :   assert (rdbk == 32'd10335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	366   :   assert (rdbk == 32'd11066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	367   :   assert (rdbk == 32'd11799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	368   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	369   :   assert (rdbk == 32'd982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	370   :   assert (rdbk == 32'd1721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	371   :   assert (rdbk == 32'd2462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	372   :   assert (rdbk == 32'd3205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	373   :   assert (rdbk == 32'd3950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	374   :   assert (rdbk == 32'd4697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	375   :   assert (rdbk == 32'd5446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	376   :   assert (rdbk == 32'd6197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	377   :   assert (rdbk == 32'd6950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	378   :   assert (rdbk == 32'd7705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	379   :   assert (rdbk == 32'd8462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	380   :   assert (rdbk == 32'd9221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	381   :   assert (rdbk == 32'd9982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	382   :   assert (rdbk == 32'd10745) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	383   :   assert (rdbk == 32'd11510) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	384   :   assert (rdbk == 32'd12277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	385   :   assert (rdbk == 32'd757) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	386   :   assert (rdbk == 32'd1528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	387   :   assert (rdbk == 32'd2301) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	388   :   assert (rdbk == 32'd3076) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	389   :   assert (rdbk == 32'd3853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	390   :   assert (rdbk == 32'd4632) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	391   :   assert (rdbk == 32'd5413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	392   :   assert (rdbk == 32'd6196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	393   :   assert (rdbk == 32'd6981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	394   :   assert (rdbk == 32'd7768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	395   :   assert (rdbk == 32'd8557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	396   :   assert (rdbk == 32'd9348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	397   :   assert (rdbk == 32'd10141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	398   :   assert (rdbk == 32'd10936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	399   :   assert (rdbk == 32'd11733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	400   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	401   :   assert (rdbk == 32'd1044) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	402   :   assert (rdbk == 32'd1847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	403   :   assert (rdbk == 32'd2652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	404   :   assert (rdbk == 32'd3459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	405   :   assert (rdbk == 32'd4268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	406   :   assert (rdbk == 32'd5079) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	407   :   assert (rdbk == 32'd5892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	408   :   assert (rdbk == 32'd6707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	409   :   assert (rdbk == 32'd7524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	410   :   assert (rdbk == 32'd8343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	411   :   assert (rdbk == 32'd9164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	412   :   assert (rdbk == 32'd9987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	413   :   assert (rdbk == 32'd10812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	414   :   assert (rdbk == 32'd11639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	415   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	416   :   assert (rdbk == 32'd1010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	417   :   assert (rdbk == 32'd1843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	418   :   assert (rdbk == 32'd2678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	419   :   assert (rdbk == 32'd3515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	420   :   assert (rdbk == 32'd4354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	421   :   assert (rdbk == 32'd5195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	422   :   assert (rdbk == 32'd6038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	423   :   assert (rdbk == 32'd6883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	424   :   assert (rdbk == 32'd7730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	425   :   assert (rdbk == 32'd8579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	426   :   assert (rdbk == 32'd9430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	427   :   assert (rdbk == 32'd10283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	428   :   assert (rdbk == 32'd11138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	429   :   assert (rdbk == 32'd11995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	430   :   assert (rdbk == 32'd565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	431   :   assert (rdbk == 32'd1426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	432   :   assert (rdbk == 32'd2289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	433   :   assert (rdbk == 32'd3154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	434   :   assert (rdbk == 32'd4021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	435   :   assert (rdbk == 32'd4890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	436   :   assert (rdbk == 32'd5761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	437   :   assert (rdbk == 32'd6634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	438   :   assert (rdbk == 32'd7509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	439   :   assert (rdbk == 32'd8386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	440   :   assert (rdbk == 32'd9265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	441   :   assert (rdbk == 32'd10146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	442   :   assert (rdbk == 32'd11029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	443   :   assert (rdbk == 32'd11914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	444   :   assert (rdbk == 32'd512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	445   :   assert (rdbk == 32'd1401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	446   :   assert (rdbk == 32'd2292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	447   :   assert (rdbk == 32'd3185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	448   :   assert (rdbk == 32'd4080) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	449   :   assert (rdbk == 32'd4977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	450   :   assert (rdbk == 32'd5876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	451   :   assert (rdbk == 32'd6777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	452   :   assert (rdbk == 32'd7680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	453   :   assert (rdbk == 32'd8585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	454   :   assert (rdbk == 32'd9492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	455   :   assert (rdbk == 32'd10401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	456   :   assert (rdbk == 32'd11312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	457   :   assert (rdbk == 32'd12225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	458   :   assert (rdbk == 32'd851) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	459   :   assert (rdbk == 32'd1768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	460   :   assert (rdbk == 32'd2687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	461   :   assert (rdbk == 32'd3608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	462   :   assert (rdbk == 32'd4531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	463   :   assert (rdbk == 32'd5456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	464   :   assert (rdbk == 32'd6383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	465   :   assert (rdbk == 32'd7312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	466   :   assert (rdbk == 32'd8243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	467   :   assert (rdbk == 32'd9176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	468   :   assert (rdbk == 32'd10111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	469   :   assert (rdbk == 32'd11048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	470   :   assert (rdbk == 32'd11987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	471   :   assert (rdbk == 32'd639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	472   :   assert (rdbk == 32'd1582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	473   :   assert (rdbk == 32'd2527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	474   :   assert (rdbk == 32'd3474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	475   :   assert (rdbk == 32'd4423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	476   :   assert (rdbk == 32'd5374) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	477   :   assert (rdbk == 32'd6327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	478   :   assert (rdbk == 32'd7282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	479   :   assert (rdbk == 32'd8239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	480   :   assert (rdbk == 32'd9198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	481   :   assert (rdbk == 32'd10159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	482   :   assert (rdbk == 32'd11122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	483   :   assert (rdbk == 32'd12087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	484   :   assert (rdbk == 32'd765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	485   :   assert (rdbk == 32'd1734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	486   :   assert (rdbk == 32'd2705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	487   :   assert (rdbk == 32'd3678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	488   :   assert (rdbk == 32'd4653) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	489   :   assert (rdbk == 32'd5630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	490   :   assert (rdbk == 32'd6609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	491   :   assert (rdbk == 32'd7590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	492   :   assert (rdbk == 32'd8573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	493   :   assert (rdbk == 32'd9558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	494   :   assert (rdbk == 32'd10545) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	495   :   assert (rdbk == 32'd11534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	496   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	497   :   assert (rdbk == 32'd1229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	498   :   assert (rdbk == 32'd2224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	499   :   assert (rdbk == 32'd3221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	500   :   assert (rdbk == 32'd4220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	501   :   assert (rdbk == 32'd5221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	502   :   assert (rdbk == 32'd6224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	503   :   assert (rdbk == 32'd7229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	504   :   assert (rdbk == 32'd8236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	505   :   assert (rdbk == 32'd9245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	506   :   assert (rdbk == 32'd10256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	507   :   assert (rdbk == 32'd11269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	508   :   assert (rdbk == 32'd12284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	509   :   assert (rdbk == 32'd1012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	510   :   assert (rdbk == 32'd2031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	511   :   assert (rdbk == 32'd3052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	512   :   assert (rdbk == 32'd4075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	513   :   assert (rdbk == 32'd5100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	514   :   assert (rdbk == 32'd6127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	515   :   assert (rdbk == 32'd7156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	516   :   assert (rdbk == 32'd8187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	517   :   assert (rdbk == 32'd9220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	518   :   assert (rdbk == 32'd10255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	519   :   assert (rdbk == 32'd11292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	520   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	521   :   assert (rdbk == 32'd1083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	522   :   assert (rdbk == 32'd2126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	523   :   assert (rdbk == 32'd3171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	524   :   assert (rdbk == 32'd4218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	525   :   assert (rdbk == 32'd5267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	526   :   assert (rdbk == 32'd6318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	527   :   assert (rdbk == 32'd7371) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	528   :   assert (rdbk == 32'd8426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	529   :   assert (rdbk == 32'd9483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	530   :   assert (rdbk == 32'd10542) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	531   :   assert (rdbk == 32'd11603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	532   :   assert (rdbk == 32'd377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	533   :   assert (rdbk == 32'd1442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	534   :   assert (rdbk == 32'd2509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	535   :   assert (rdbk == 32'd3578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	536   :   assert (rdbk == 32'd4649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	537   :   assert (rdbk == 32'd5722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	538   :   assert (rdbk == 32'd6797) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	539   :   assert (rdbk == 32'd7874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	540   :   assert (rdbk == 32'd8953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	541   :   assert (rdbk == 32'd10034) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	542   :   assert (rdbk == 32'd11117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	543   :   assert (rdbk == 32'd12202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	544   :   assert (rdbk == 32'd1000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	545   :   assert (rdbk == 32'd2089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	546   :   assert (rdbk == 32'd3180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	547   :   assert (rdbk == 32'd4273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	548   :   assert (rdbk == 32'd5368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	549   :   assert (rdbk == 32'd6465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	550   :   assert (rdbk == 32'd7564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	551   :   assert (rdbk == 32'd8665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	552   :   assert (rdbk == 32'd9768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	553   :   assert (rdbk == 32'd10873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	554   :   assert (rdbk == 32'd11980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	555   :   assert (rdbk == 32'd800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	556   :   assert (rdbk == 32'd1911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	557   :   assert (rdbk == 32'd3024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	558   :   assert (rdbk == 32'd4139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	559   :   assert (rdbk == 32'd5256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	560   :   assert (rdbk == 32'd6375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	561   :   assert (rdbk == 32'd7496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	562   :   assert (rdbk == 32'd8619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	563   :   assert (rdbk == 32'd9744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	564   :   assert (rdbk == 32'd10871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	565   :   assert (rdbk == 32'd12000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	566   :   assert (rdbk == 32'd842) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	567   :   assert (rdbk == 32'd1975) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	568   :   assert (rdbk == 32'd3110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	569   :   assert (rdbk == 32'd4247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	570   :   assert (rdbk == 32'd5386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	571   :   assert (rdbk == 32'd6527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	572   :   assert (rdbk == 32'd7670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	573   :   assert (rdbk == 32'd8815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	574   :   assert (rdbk == 32'd9962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	575   :   assert (rdbk == 32'd11111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	576   :   assert (rdbk == 32'd12262) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	577   :   assert (rdbk == 32'd1126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	578   :   assert (rdbk == 32'd2281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	579   :   assert (rdbk == 32'd3438) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	580   :   assert (rdbk == 32'd4597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	581   :   assert (rdbk == 32'd5758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	582   :   assert (rdbk == 32'd6921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	583   :   assert (rdbk == 32'd8086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	584   :   assert (rdbk == 32'd9253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	585   :   assert (rdbk == 32'd10422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	586   :   assert (rdbk == 32'd11593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	587   :   assert (rdbk == 32'd477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	588   :   assert (rdbk == 32'd1652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	589   :   assert (rdbk == 32'd2829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	590   :   assert (rdbk == 32'd4008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	591   :   assert (rdbk == 32'd5189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	592   :   assert (rdbk == 32'd6372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	593   :   assert (rdbk == 32'd7557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	594   :   assert (rdbk == 32'd8744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	595   :   assert (rdbk == 32'd9933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	596   :   assert (rdbk == 32'd11124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	597   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	598   :   assert (rdbk == 32'd1223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	599   :   assert (rdbk == 32'd2420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	600   :   assert (rdbk == 32'd3619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	601   :   assert (rdbk == 32'd4820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	602   :   assert (rdbk == 32'd6023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	603   :   assert (rdbk == 32'd7228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	604   :   assert (rdbk == 32'd8435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	605   :   assert (rdbk == 32'd9644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	606   :   assert (rdbk == 32'd10855) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	607   :   assert (rdbk == 32'd12068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	608   :   assert (rdbk == 32'd994) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	609   :   assert (rdbk == 32'd2211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	610   :   assert (rdbk == 32'd3430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	611   :   assert (rdbk == 32'd4651) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	612   :   assert (rdbk == 32'd5874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	613   :   assert (rdbk == 32'd7099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	614   :   assert (rdbk == 32'd8326) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	615   :   assert (rdbk == 32'd9555) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	616   :   assert (rdbk == 32'd10786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	617   :   assert (rdbk == 32'd12019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	618   :   assert (rdbk == 32'd965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	619   :   assert (rdbk == 32'd2202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	620   :   assert (rdbk == 32'd3441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	621   :   assert (rdbk == 32'd4682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	622   :   assert (rdbk == 32'd5925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	623   :   assert (rdbk == 32'd7170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	624   :   assert (rdbk == 32'd8417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	625   :   assert (rdbk == 32'd9666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	626   :   assert (rdbk == 32'd10917) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	627   :   assert (rdbk == 32'd12170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	628   :   assert (rdbk == 32'd1136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	629   :   assert (rdbk == 32'd2393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	630   :   assert (rdbk == 32'd3652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	631   :   assert (rdbk == 32'd4913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	632   :   assert (rdbk == 32'd6176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	633   :   assert (rdbk == 32'd7441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	634   :   assert (rdbk == 32'd8708) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	635   :   assert (rdbk == 32'd9977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	636   :   assert (rdbk == 32'd11248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	637   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	638   :   assert (rdbk == 32'd1507) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	639   :   assert (rdbk == 32'd2784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	640   :   assert (rdbk == 32'd4063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	641   :   assert (rdbk == 32'd5344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	642   :   assert (rdbk == 32'd6627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	643   :   assert (rdbk == 32'd7912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	644   :   assert (rdbk == 32'd9199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	645   :   assert (rdbk == 32'd10488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	646   :   assert (rdbk == 32'd11779) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	647   :   assert (rdbk == 32'd783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	648   :   assert (rdbk == 32'd2078) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	649   :   assert (rdbk == 32'd3375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	650   :   assert (rdbk == 32'd4674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	651   :   assert (rdbk == 32'd5975) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	652   :   assert (rdbk == 32'd7278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	653   :   assert (rdbk == 32'd8583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	654   :   assert (rdbk == 32'd9890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	655   :   assert (rdbk == 32'd11199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	656   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	657   :   assert (rdbk == 32'd1534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	658   :   assert (rdbk == 32'd2849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	659   :   assert (rdbk == 32'd4166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	660   :   assert (rdbk == 32'd5485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	661   :   assert (rdbk == 32'd6806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	662   :   assert (rdbk == 32'd8129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	663   :   assert (rdbk == 32'd9454) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	664   :   assert (rdbk == 32'd10781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	665   :   assert (rdbk == 32'd12110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	666   :   assert (rdbk == 32'd1152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	667   :   assert (rdbk == 32'd2485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	668   :   assert (rdbk == 32'd3820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	669   :   assert (rdbk == 32'd5157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	670   :   assert (rdbk == 32'd6496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	671   :   assert (rdbk == 32'd7837) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	672   :   assert (rdbk == 32'd9180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	673   :   assert (rdbk == 32'd10525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	674   :   assert (rdbk == 32'd11872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	675   :   assert (rdbk == 32'd932) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	676   :   assert (rdbk == 32'd2283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	677   :   assert (rdbk == 32'd3636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	678   :   assert (rdbk == 32'd4991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	679   :   assert (rdbk == 32'd6348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	680   :   assert (rdbk == 32'd7707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	681   :   assert (rdbk == 32'd9068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	682   :   assert (rdbk == 32'd10431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	683   :   assert (rdbk == 32'd11796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	684   :   assert (rdbk == 32'd874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	685   :   assert (rdbk == 32'd2243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	686   :   assert (rdbk == 32'd3614) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	687   :   assert (rdbk == 32'd4987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	688   :   assert (rdbk == 32'd6362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	689   :   assert (rdbk == 32'd7739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	690   :   assert (rdbk == 32'd9118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	691   :   assert (rdbk == 32'd10499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	692   :   assert (rdbk == 32'd11882) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	693   :   assert (rdbk == 32'd978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	694   :   assert (rdbk == 32'd2365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	695   :   assert (rdbk == 32'd3754) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	696   :   assert (rdbk == 32'd5145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	697   :   assert (rdbk == 32'd6538) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	698   :   assert (rdbk == 32'd7933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	699   :   assert (rdbk == 32'd9330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	700   :   assert (rdbk == 32'd10729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	701   :   assert (rdbk == 32'd12130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	702   :   assert (rdbk == 32'd1244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	703   :   assert (rdbk == 32'd2649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	704   :   assert (rdbk == 32'd4056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	705   :   assert (rdbk == 32'd5465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	706   :   assert (rdbk == 32'd6876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	707   :   assert (rdbk == 32'd8289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	708   :   assert (rdbk == 32'd9704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	709   :   assert (rdbk == 32'd11121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	710   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	711   :   assert (rdbk == 32'd1672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	712   :   assert (rdbk == 32'd3095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	713   :   assert (rdbk == 32'd4520) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	714   :   assert (rdbk == 32'd5947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	715   :   assert (rdbk == 32'd7376) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	716   :   assert (rdbk == 32'd8807) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	717   :   assert (rdbk == 32'd10240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	718   :   assert (rdbk == 32'd11675) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	719   :   assert (rdbk == 32'd823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	720   :   assert (rdbk == 32'd2262) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	721   :   assert (rdbk == 32'd3703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	722   :   assert (rdbk == 32'd5146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	723   :   assert (rdbk == 32'd6591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	724   :   assert (rdbk == 32'd8038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	725   :   assert (rdbk == 32'd9487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	726   :   assert (rdbk == 32'd10938) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	727   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	728   :   assert (rdbk == 32'd1557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	729   :   assert (rdbk == 32'd3014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	730   :   assert (rdbk == 32'd4473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	731   :   assert (rdbk == 32'd5934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	732   :   assert (rdbk == 32'd7397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	733   :   assert (rdbk == 32'd8862) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	734   :   assert (rdbk == 32'd10329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	735   :   assert (rdbk == 32'd11798) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	736   :   assert (rdbk == 32'd980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	737   :   assert (rdbk == 32'd2453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	738   :   assert (rdbk == 32'd3928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	739   :   assert (rdbk == 32'd5405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	740   :   assert (rdbk == 32'd6884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	741   :   assert (rdbk == 32'd8365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	742   :   assert (rdbk == 32'd9848) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	743   :   assert (rdbk == 32'd11333) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	744   :   assert (rdbk == 32'd531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	745   :   assert (rdbk == 32'd2020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	746   :   assert (rdbk == 32'd3511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	747   :   assert (rdbk == 32'd5004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	748   :   assert (rdbk == 32'd6499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	749   :   assert (rdbk == 32'd7996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	750   :   assert (rdbk == 32'd9495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	751   :   assert (rdbk == 32'd10996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	752   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	753   :   assert (rdbk == 32'd1715) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	754   :   assert (rdbk == 32'd3222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	755   :   assert (rdbk == 32'd4731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	756   :   assert (rdbk == 32'd6242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	757   :   assert (rdbk == 32'd7755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	758   :   assert (rdbk == 32'd9270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	759   :   assert (rdbk == 32'd10787) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	760   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	761   :   assert (rdbk == 32'd1538) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	762   :   assert (rdbk == 32'd3061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	763   :   assert (rdbk == 32'd4586) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	764   :   assert (rdbk == 32'd6113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	765   :   assert (rdbk == 32'd7642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	766   :   assert (rdbk == 32'd9173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	767   :   assert (rdbk == 32'd10706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	768   :   assert (rdbk == 32'd12241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	769   :   assert (rdbk == 32'd1489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	770   :   assert (rdbk == 32'd3028) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	771   :   assert (rdbk == 32'd4569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	772   :   assert (rdbk == 32'd6112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	773   :   assert (rdbk == 32'd7657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	774   :   assert (rdbk == 32'd9204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	775   :   assert (rdbk == 32'd10753) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	776   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	777   :   assert (rdbk == 32'd1568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	778   :   assert (rdbk == 32'd3123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	779   :   assert (rdbk == 32'd4680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	780   :   assert (rdbk == 32'd6239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	781   :   assert (rdbk == 32'd7800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	782   :   assert (rdbk == 32'd9363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	783   :   assert (rdbk == 32'd10928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	784   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	785   :   assert (rdbk == 32'd1775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	786   :   assert (rdbk == 32'd3346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	787   :   assert (rdbk == 32'd4919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	788   :   assert (rdbk == 32'd6494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	789   :   assert (rdbk == 32'd8071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	790   :   assert (rdbk == 32'd9650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	791   :   assert (rdbk == 32'd11231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	792   :   assert (rdbk == 32'd525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	793   :   assert (rdbk == 32'd2110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	794   :   assert (rdbk == 32'd3697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	795   :   assert (rdbk == 32'd5286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	796   :   assert (rdbk == 32'd6877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	797   :   assert (rdbk == 32'd8470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	798   :   assert (rdbk == 32'd10065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	799   :   assert (rdbk == 32'd11662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	800   :   assert (rdbk == 32'd972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	801   :   assert (rdbk == 32'd2573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	802   :   assert (rdbk == 32'd4176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	803   :   assert (rdbk == 32'd5781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	804   :   assert (rdbk == 32'd7388) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	805   :   assert (rdbk == 32'd8997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	806   :   assert (rdbk == 32'd10608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	807   :   assert (rdbk == 32'd12221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	808   :   assert (rdbk == 32'd1547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	809   :   assert (rdbk == 32'd3164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	810   :   assert (rdbk == 32'd4783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	811   :   assert (rdbk == 32'd6404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	812   :   assert (rdbk == 32'd8027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	813   :   assert (rdbk == 32'd9652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	814   :   assert (rdbk == 32'd11279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	815   :   assert (rdbk == 32'd619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	816   :   assert (rdbk == 32'd2250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	817   :   assert (rdbk == 32'd3883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	818   :   assert (rdbk == 32'd5518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	819   :   assert (rdbk == 32'd7155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	820   :   assert (rdbk == 32'd8794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	821   :   assert (rdbk == 32'd10435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	822   :   assert (rdbk == 32'd12078) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	823   :   assert (rdbk == 32'd1434) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	824   :   assert (rdbk == 32'd3081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	825   :   assert (rdbk == 32'd4730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	826   :   assert (rdbk == 32'd6381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	827   :   assert (rdbk == 32'd8034) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	828   :   assert (rdbk == 32'd9689) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	829   :   assert (rdbk == 32'd11346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	830   :   assert (rdbk == 32'd716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	831   :   assert (rdbk == 32'd2377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	832   :   assert (rdbk == 32'd4040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	833   :   assert (rdbk == 32'd5705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	834   :   assert (rdbk == 32'd7372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	835   :   assert (rdbk == 32'd9041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	836   :   assert (rdbk == 32'd10712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	837   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	838   :   assert (rdbk == 32'd1771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	839   :   assert (rdbk == 32'd3448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	840   :   assert (rdbk == 32'd5127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	841   :   assert (rdbk == 32'd6808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	842   :   assert (rdbk == 32'd8491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	843   :   assert (rdbk == 32'd10176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	844   :   assert (rdbk == 32'd11863) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	845   :   assert (rdbk == 32'd1263) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	846   :   assert (rdbk == 32'd2954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	847   :   assert (rdbk == 32'd4647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	848   :   assert (rdbk == 32'd6342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	849   :   assert (rdbk == 32'd8039) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	850   :   assert (rdbk == 32'd9738) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	851   :   assert (rdbk == 32'd11439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	852   :   assert (rdbk == 32'd853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	853   :   assert (rdbk == 32'd2558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	854   :   assert (rdbk == 32'd4265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	855   :   assert (rdbk == 32'd5974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	856   :   assert (rdbk == 32'd7685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	857   :   assert (rdbk == 32'd9398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	858   :   assert (rdbk == 32'd11113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	859   :   assert (rdbk == 32'd541) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	860   :   assert (rdbk == 32'd2260) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	861   :   assert (rdbk == 32'd3981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	862   :   assert (rdbk == 32'd5704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	863   :   assert (rdbk == 32'd7429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	864   :   assert (rdbk == 32'd9156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	865   :   assert (rdbk == 32'd10885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	866   :   assert (rdbk == 32'd327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	867   :   assert (rdbk == 32'd2060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	868   :   assert (rdbk == 32'd3795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	869   :   assert (rdbk == 32'd5532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	870   :   assert (rdbk == 32'd7271) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	871   :   assert (rdbk == 32'd9012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	872   :   assert (rdbk == 32'd10755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	873   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	874   :   assert (rdbk == 32'd1958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	875   :   assert (rdbk == 32'd3707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	876   :   assert (rdbk == 32'd5458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	877   :   assert (rdbk == 32'd7211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	878   :   assert (rdbk == 32'd8966) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	879   :   assert (rdbk == 32'd10723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	880   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	881   :   assert (rdbk == 32'd1954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	882   :   assert (rdbk == 32'd3717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	883   :   assert (rdbk == 32'd5482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	884   :   assert (rdbk == 32'd7249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	885   :   assert (rdbk == 32'd9018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	886   :   assert (rdbk == 32'd10789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	887   :   assert (rdbk == 32'd273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	888   :   assert (rdbk == 32'd2048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	889   :   assert (rdbk == 32'd3825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	890   :   assert (rdbk == 32'd5604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	891   :   assert (rdbk == 32'd7385) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	892   :   assert (rdbk == 32'd9168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	893   :   assert (rdbk == 32'd10953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	894   :   assert (rdbk == 32'd451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	895   :   assert (rdbk == 32'd2240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	896   :   assert (rdbk == 32'd4031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	897   :   assert (rdbk == 32'd5824) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	898   :   assert (rdbk == 32'd7619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	899   :   assert (rdbk == 32'd9416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	900   :   assert (rdbk == 32'd11215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	901   :   assert (rdbk == 32'd727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	902   :   assert (rdbk == 32'd2530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	903   :   assert (rdbk == 32'd4335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	904   :   assert (rdbk == 32'd6142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	905   :   assert (rdbk == 32'd7951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	906   :   assert (rdbk == 32'd9762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	907   :   assert (rdbk == 32'd11575) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	908   :   assert (rdbk == 32'd1101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	909   :   assert (rdbk == 32'd2918) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	910   :   assert (rdbk == 32'd4737) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	911   :   assert (rdbk == 32'd6558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	912   :   assert (rdbk == 32'd8381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	913   :   assert (rdbk == 32'd10206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	914   :   assert (rdbk == 32'd12033) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	915   :   assert (rdbk == 32'd1573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	916   :   assert (rdbk == 32'd3404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	917   :   assert (rdbk == 32'd5237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	918   :   assert (rdbk == 32'd7072) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	919   :   assert (rdbk == 32'd8909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	920   :   assert (rdbk == 32'd10748) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	921   :   assert (rdbk == 32'd300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	922   :   assert (rdbk == 32'd2143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	923   :   assert (rdbk == 32'd3988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	924   :   assert (rdbk == 32'd5835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	925   :   assert (rdbk == 32'd7684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	926   :   assert (rdbk == 32'd9535) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	927   :   assert (rdbk == 32'd11388) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	928   :   assert (rdbk == 32'd954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	929   :   assert (rdbk == 32'd2811) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	930   :   assert (rdbk == 32'd4670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	931   :   assert (rdbk == 32'd6531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	932   :   assert (rdbk == 32'd8394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	933   :   assert (rdbk == 32'd10259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	934   :   assert (rdbk == 32'd12126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	935   :   assert (rdbk == 32'd1706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	936   :   assert (rdbk == 32'd3577) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	937   :   assert (rdbk == 32'd5450) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	938   :   assert (rdbk == 32'd7325) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	939   :   assert (rdbk == 32'd9202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	940   :   assert (rdbk == 32'd11081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	941   :   assert (rdbk == 32'd673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	942   :   assert (rdbk == 32'd2556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	943   :   assert (rdbk == 32'd4441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	944   :   assert (rdbk == 32'd6328) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	945   :   assert (rdbk == 32'd8217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	946   :   assert (rdbk == 32'd10108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	947   :   assert (rdbk == 32'd12001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	948   :   assert (rdbk == 32'd1607) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	949   :   assert (rdbk == 32'd3504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	950   :   assert (rdbk == 32'd5403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	951   :   assert (rdbk == 32'd7304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	952   :   assert (rdbk == 32'd9207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	953   :   assert (rdbk == 32'd11112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	954   :   assert (rdbk == 32'd730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	955   :   assert (rdbk == 32'd2639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	956   :   assert (rdbk == 32'd4550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	957   :   assert (rdbk == 32'd6463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	958   :   assert (rdbk == 32'd8378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	959   :   assert (rdbk == 32'd10295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	960   :   assert (rdbk == 32'd12214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	961   :   assert (rdbk == 32'd1846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	962   :   assert (rdbk == 32'd3769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	963   :   assert (rdbk == 32'd5694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	964   :   assert (rdbk == 32'd7621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	965   :   assert (rdbk == 32'd9550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	966   :   assert (rdbk == 32'd11481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	967   :   assert (rdbk == 32'd1125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	968   :   assert (rdbk == 32'd3060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	969   :   assert (rdbk == 32'd4997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	970   :   assert (rdbk == 32'd6936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	971   :   assert (rdbk == 32'd8877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	972   :   assert (rdbk == 32'd10820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	973   :   assert (rdbk == 32'd476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	974   :   assert (rdbk == 32'd2423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	975   :   assert (rdbk == 32'd4372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	976   :   assert (rdbk == 32'd6323) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	977   :   assert (rdbk == 32'd8276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	978   :   assert (rdbk == 32'd10231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	979   :   assert (rdbk == 32'd12188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	980   :   assert (rdbk == 32'd1858) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	981   :   assert (rdbk == 32'd3819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	982   :   assert (rdbk == 32'd5782) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	983   :   assert (rdbk == 32'd7747) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	984   :   assert (rdbk == 32'd9714) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	985   :   assert (rdbk == 32'd11683) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	986   :   assert (rdbk == 32'd1365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	987   :   assert (rdbk == 32'd3338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	988   :   assert (rdbk == 32'd5313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	989   :   assert (rdbk == 32'd7290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	990   :   assert (rdbk == 32'd9269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	991   :   assert (rdbk == 32'd11250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	992   :   assert (rdbk == 32'd944) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	993   :   assert (rdbk == 32'd2929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	994   :   assert (rdbk == 32'd4916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	995   :   assert (rdbk == 32'd6905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	996   :   assert (rdbk == 32'd8896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	997   :   assert (rdbk == 32'd10889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	998   :   assert (rdbk == 32'd595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	999   :   assert (rdbk == 32'd2592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1000   :   assert (rdbk == 32'd4591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1001   :   assert (rdbk == 32'd6592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1002   :   assert (rdbk == 32'd8595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1003   :   assert (rdbk == 32'd10600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1004   :   assert (rdbk == 32'd318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1005   :   assert (rdbk == 32'd2327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1006   :   assert (rdbk == 32'd4338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1007   :   assert (rdbk == 32'd6351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1008   :   assert (rdbk == 32'd8366) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1009   :   assert (rdbk == 32'd10383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1010   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1011   :   assert (rdbk == 32'd2134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1012   :   assert (rdbk == 32'd4157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1013   :   assert (rdbk == 32'd6182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1014   :   assert (rdbk == 32'd8209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1015   :   assert (rdbk == 32'd10238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1016   :   assert (rdbk == 32'd12269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1017   :   assert (rdbk == 32'd2013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1018   :   assert (rdbk == 32'd4048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1019   :   assert (rdbk == 32'd6085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1020   :   assert (rdbk == 32'd8124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1021   :   assert (rdbk == 32'd10165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1022   :   assert (rdbk == 32'd12208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1023   :   assert (rdbk == 32'd1964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
    endcase
end

