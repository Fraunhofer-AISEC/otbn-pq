// Copyright Copyright Fraunhofer Institute for Applied and Integrated Security (AISEC).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

$fwrite(f,"----------------------------------------------------------------\n");   
$fwrite(f,"-- Falcon-1024 - Singature Verification Test \n");
$fwrite(f,"----------------------------------------------------------------\n");   
     
// Write IMEM from File
write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq_falcon1024-valid.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- IMEM\n");
// Read IMEM  
for (int i=0 ; i<129 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end     

 // Write DMEM from File
write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq_falcon1024-valid.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- DMEM\n");
// Read DMEM  
for (int i=0 ; i<16 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end   
	   
$fwrite(f,"----------------------------------------------------------------\n");   

// Set Instruction Counter to zero (optional)
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );

// Start Programm in IMEM
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(CmdExecute), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
cc_start = cc;
// Poll on Status Register until Programm is finished
rdbk = '1;
while (rdbk != '0) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
end 

// Measure CC
cc_stop = cc; 
cc_count_falcon1024_1 = cc_stop - cc_start;        
       
// Read DMEM  
for (int i=0 ; i<1024 ; i++) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+448+4096*3), .tl_o(tl_o), .tl_i(tl_i_d) );
    
    case(i)
	0   :   assert (rdbk == 32'h0000004c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1   :   assert (rdbk == 32'hffffffdf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2   :   assert (rdbk == 32'h0000004d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3   :   assert (rdbk == 32'hffffffa1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4   :   assert (rdbk == 32'hfffffecd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	5   :   assert (rdbk == 32'hffffff9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	6   :   assert (rdbk == 32'h000000a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	7   :   assert (rdbk == 32'h00000050) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	8   :   assert (rdbk == 32'hffffff90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	9   :   assert (rdbk == 32'h00000088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	10   :   assert (rdbk == 32'hffffff66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	11   :   assert (rdbk == 32'hffffff75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	12   :   assert (rdbk == 32'hffffff8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	13   :   assert (rdbk == 32'h000000d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	14   :   assert (rdbk == 32'hffffffd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	15   :   assert (rdbk == 32'h000000ae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	16   :   assert (rdbk == 32'hffffffd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	17   :   assert (rdbk == 32'hffffff6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	18   :   assert (rdbk == 32'h0000001e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	19   :   assert (rdbk == 32'hffffff2b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	20   :   assert (rdbk == 32'hffffff84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	21   :   assert (rdbk == 32'h000001cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	22   :   assert (rdbk == 32'hfffffed6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	23   :   assert (rdbk == 32'hffffffec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	24   :   assert (rdbk == 32'hfffffeb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	25   :   assert (rdbk == 32'h00000011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	26   :   assert (rdbk == 32'h0000005d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	27   :   assert (rdbk == 32'h00000013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	28   :   assert (rdbk == 32'hfffffff8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	29   :   assert (rdbk == 32'h0000006a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	30   :   assert (rdbk == 32'hffffffbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	31   :   assert (rdbk == 32'hffffff95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	32   :   assert (rdbk == 32'h0000001c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	33   :   assert (rdbk == 32'h000000e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	34   :   assert (rdbk == 32'hffffffe3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	35   :   assert (rdbk == 32'hffffff6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	36   :   assert (rdbk == 32'hffffff5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	37   :   assert (rdbk == 32'h000001ef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	38   :   assert (rdbk == 32'h000000ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	39   :   assert (rdbk == 32'h00000085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	40   :   assert (rdbk == 32'hffffff6b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	41   :   assert (rdbk == 32'h00000000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	42   :   assert (rdbk == 32'h0000004d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	43   :   assert (rdbk == 32'h00000108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	44   :   assert (rdbk == 32'hfffffff7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	45   :   assert (rdbk == 32'h0000003f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	46   :   assert (rdbk == 32'hffffffea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	47   :   assert (rdbk == 32'h00000001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	48   :   assert (rdbk == 32'h0000001c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	49   :   assert (rdbk == 32'hffffff8d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	50   :   assert (rdbk == 32'hffffff7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	51   :   assert (rdbk == 32'hffffffce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	52   :   assert (rdbk == 32'hffffff71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	53   :   assert (rdbk == 32'hffffffbb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	54   :   assert (rdbk == 32'h00000010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	55   :   assert (rdbk == 32'hffffffcf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	56   :   assert (rdbk == 32'hffffff9e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	57   :   assert (rdbk == 32'hffffffb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	58   :   assert (rdbk == 32'hffffffa3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	59   :   assert (rdbk == 32'h00000100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	60   :   assert (rdbk == 32'hffffffed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	61   :   assert (rdbk == 32'hffffffde) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	62   :   assert (rdbk == 32'h0000003b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	63   :   assert (rdbk == 32'h0000000c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	64   :   assert (rdbk == 32'hffffffcf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	65   :   assert (rdbk == 32'hffffffe2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	66   :   assert (rdbk == 32'hfffffefb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	67   :   assert (rdbk == 32'hffffffb4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	68   :   assert (rdbk == 32'h000000d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	69   :   assert (rdbk == 32'h00000054) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	70   :   assert (rdbk == 32'h000000bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	71   :   assert (rdbk == 32'h0000008b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	72   :   assert (rdbk == 32'h0000004a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	73   :   assert (rdbk == 32'h000000ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	74   :   assert (rdbk == 32'hfffffec5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	75   :   assert (rdbk == 32'h000000fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	76   :   assert (rdbk == 32'hffffffbe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	77   :   assert (rdbk == 32'h00000050) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	78   :   assert (rdbk == 32'h00000037) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	79   :   assert (rdbk == 32'h000000c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	80   :   assert (rdbk == 32'h0000003a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	81   :   assert (rdbk == 32'h0000000f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	82   :   assert (rdbk == 32'hffffff8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	83   :   assert (rdbk == 32'hffffff6d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	84   :   assert (rdbk == 32'h00000014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	85   :   assert (rdbk == 32'h0000006c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	86   :   assert (rdbk == 32'h0000014b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	87   :   assert (rdbk == 32'hffffffdc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	88   :   assert (rdbk == 32'hffffff8d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	89   :   assert (rdbk == 32'h00000123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	90   :   assert (rdbk == 32'hffffffc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	91   :   assert (rdbk == 32'h00000097) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	92   :   assert (rdbk == 32'hffffff8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	93   :   assert (rdbk == 32'hffffff45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	94   :   assert (rdbk == 32'hffffff84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	95   :   assert (rdbk == 32'h00000066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	96   :   assert (rdbk == 32'h00000069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	97   :   assert (rdbk == 32'h000000c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	98   :   assert (rdbk == 32'h00000068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	99   :   assert (rdbk == 32'hffffff68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	100   :   assert (rdbk == 32'h00000081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	101   :   assert (rdbk == 32'h000000ec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	102   :   assert (rdbk == 32'h0000002a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	103   :   assert (rdbk == 32'hffffff97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	104   :   assert (rdbk == 32'hffffffa0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	105   :   assert (rdbk == 32'h0000003d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	106   :   assert (rdbk == 32'h00000069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	107   :   assert (rdbk == 32'h0000003a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	108   :   assert (rdbk == 32'h0000000d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	109   :   assert (rdbk == 32'hfffffffd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	110   :   assert (rdbk == 32'h0000003f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	111   :   assert (rdbk == 32'h000000a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	112   :   assert (rdbk == 32'hffffff12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	113   :   assert (rdbk == 32'h00000142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	114   :   assert (rdbk == 32'h00000063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	115   :   assert (rdbk == 32'h00000012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	116   :   assert (rdbk == 32'h00000000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	117   :   assert (rdbk == 32'hffffff3b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	118   :   assert (rdbk == 32'h000000b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	119   :   assert (rdbk == 32'hffffff2b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	120   :   assert (rdbk == 32'h00000099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	121   :   assert (rdbk == 32'hffffffe1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	122   :   assert (rdbk == 32'h0000010f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	123   :   assert (rdbk == 32'hffffff89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	124   :   assert (rdbk == 32'h000000a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	125   :   assert (rdbk == 32'hfffffe7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	126   :   assert (rdbk == 32'hffffff7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	127   :   assert (rdbk == 32'hffffff12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	128   :   assert (rdbk == 32'h0000006a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	129   :   assert (rdbk == 32'hffffffcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	130   :   assert (rdbk == 32'h0000008a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	131   :   assert (rdbk == 32'h0000004c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	132   :   assert (rdbk == 32'hffffff33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	133   :   assert (rdbk == 32'hffffff40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	134   :   assert (rdbk == 32'hffffffb0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	135   :   assert (rdbk == 32'hffffffb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	136   :   assert (rdbk == 32'h00000092) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	137   :   assert (rdbk == 32'h0000002a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	138   :   assert (rdbk == 32'h00000018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	139   :   assert (rdbk == 32'h000000d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	140   :   assert (rdbk == 32'hffffffb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	141   :   assert (rdbk == 32'h0000003a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	142   :   assert (rdbk == 32'hffffff57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	143   :   assert (rdbk == 32'hfffffef0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	144   :   assert (rdbk == 32'hffffffed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	145   :   assert (rdbk == 32'h0000007a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	146   :   assert (rdbk == 32'hfffffef7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	147   :   assert (rdbk == 32'h000000ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	148   :   assert (rdbk == 32'h00000055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	149   :   assert (rdbk == 32'hffffff0c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	150   :   assert (rdbk == 32'hfffffe8c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	151   :   assert (rdbk == 32'h00000032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	152   :   assert (rdbk == 32'h0000005c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	153   :   assert (rdbk == 32'h00000103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	154   :   assert (rdbk == 32'hffffffca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	155   :   assert (rdbk == 32'h000001f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	156   :   assert (rdbk == 32'h00000037) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	157   :   assert (rdbk == 32'hffffffe4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	158   :   assert (rdbk == 32'hffffffa9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	159   :   assert (rdbk == 32'h000000b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	160   :   assert (rdbk == 32'h00000072) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	161   :   assert (rdbk == 32'h0000002e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	162   :   assert (rdbk == 32'hffffffde) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	163   :   assert (rdbk == 32'h0000004d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	164   :   assert (rdbk == 32'hffffff41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	165   :   assert (rdbk == 32'h0000009a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	166   :   assert (rdbk == 32'hffffff3f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	167   :   assert (rdbk == 32'hffffff13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	168   :   assert (rdbk == 32'hffffffbc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	169   :   assert (rdbk == 32'h0000001b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	170   :   assert (rdbk == 32'hffffffb0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	171   :   assert (rdbk == 32'hffffff4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	172   :   assert (rdbk == 32'h00000091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	173   :   assert (rdbk == 32'h00000077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	174   :   assert (rdbk == 32'hffffff69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	175   :   assert (rdbk == 32'h00000047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	176   :   assert (rdbk == 32'h0000002f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	177   :   assert (rdbk == 32'h00000015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	178   :   assert (rdbk == 32'hfffffea5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	179   :   assert (rdbk == 32'h00000009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	180   :   assert (rdbk == 32'h0000001c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	181   :   assert (rdbk == 32'h0000004a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	182   :   assert (rdbk == 32'hfffffff1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	183   :   assert (rdbk == 32'hffffff87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	184   :   assert (rdbk == 32'hfffffe5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	185   :   assert (rdbk == 32'hfffffffc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	186   :   assert (rdbk == 32'hfffffffe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	187   :   assert (rdbk == 32'h0000005b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	188   :   assert (rdbk == 32'h00000166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	189   :   assert (rdbk == 32'hffffff70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	190   :   assert (rdbk == 32'hfffffec7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	191   :   assert (rdbk == 32'h0000010b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	192   :   assert (rdbk == 32'h0000004c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	193   :   assert (rdbk == 32'hffffff56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	194   :   assert (rdbk == 32'hffffffc0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	195   :   assert (rdbk == 32'h00000181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	196   :   assert (rdbk == 32'hffffff73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	197   :   assert (rdbk == 32'hffffff88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	198   :   assert (rdbk == 32'h0000013b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	199   :   assert (rdbk == 32'hffffff60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	200   :   assert (rdbk == 32'hffffffb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	201   :   assert (rdbk == 32'h0000000b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	202   :   assert (rdbk == 32'h000000e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	203   :   assert (rdbk == 32'h00000012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	204   :   assert (rdbk == 32'hffffff60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	205   :   assert (rdbk == 32'h000000bf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	206   :   assert (rdbk == 32'hfffffff8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	207   :   assert (rdbk == 32'hffffffdc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	208   :   assert (rdbk == 32'hffffffb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	209   :   assert (rdbk == 32'h00000078) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	210   :   assert (rdbk == 32'h000000e6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	211   :   assert (rdbk == 32'hffffffd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	212   :   assert (rdbk == 32'h000000a4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	213   :   assert (rdbk == 32'h00000079) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	214   :   assert (rdbk == 32'h000000e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	215   :   assert (rdbk == 32'hffffffdd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	216   :   assert (rdbk == 32'hffffffb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	217   :   assert (rdbk == 32'h00000143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	218   :   assert (rdbk == 32'h00000047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	219   :   assert (rdbk == 32'hffffff9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	220   :   assert (rdbk == 32'hffffff63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	221   :   assert (rdbk == 32'h0000010e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	222   :   assert (rdbk == 32'h00000073) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	223   :   assert (rdbk == 32'hffffffa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	224   :   assert (rdbk == 32'hffffffab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	225   :   assert (rdbk == 32'hffffffaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	226   :   assert (rdbk == 32'h00000061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	227   :   assert (rdbk == 32'h000000b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	228   :   assert (rdbk == 32'h00000031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	229   :   assert (rdbk == 32'hffffff6b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	230   :   assert (rdbk == 32'hffffffd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	231   :   assert (rdbk == 32'h00000096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	232   :   assert (rdbk == 32'hffffff83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	233   :   assert (rdbk == 32'h00000051) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	234   :   assert (rdbk == 32'hffffff4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	235   :   assert (rdbk == 32'hfffffec6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	236   :   assert (rdbk == 32'hffffffc5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	237   :   assert (rdbk == 32'hffffffc7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	238   :   assert (rdbk == 32'h0000005d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	239   :   assert (rdbk == 32'h0000008d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	240   :   assert (rdbk == 32'hffffffa1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	241   :   assert (rdbk == 32'h000000f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	242   :   assert (rdbk == 32'h00000025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	243   :   assert (rdbk == 32'h000000c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	244   :   assert (rdbk == 32'hffffffaf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	245   :   assert (rdbk == 32'h00000090) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	246   :   assert (rdbk == 32'hffffff24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	247   :   assert (rdbk == 32'h00000122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	248   :   assert (rdbk == 32'h000000fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	249   :   assert (rdbk == 32'hffffffbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	250   :   assert (rdbk == 32'hffffffdb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	251   :   assert (rdbk == 32'h000000c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	252   :   assert (rdbk == 32'h0000003b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	253   :   assert (rdbk == 32'hfffffef0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	254   :   assert (rdbk == 32'hfffffe45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	255   :   assert (rdbk == 32'h000000c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	256   :   assert (rdbk == 32'h0000001a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	257   :   assert (rdbk == 32'hffffffc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	258   :   assert (rdbk == 32'hfffffe86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	259   :   assert (rdbk == 32'hffffffe0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	260   :   assert (rdbk == 32'h000000b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	261   :   assert (rdbk == 32'h000000e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	262   :   assert (rdbk == 32'hffffffd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	263   :   assert (rdbk == 32'hffffff5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	264   :   assert (rdbk == 32'hffffff99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	265   :   assert (rdbk == 32'h000000e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	266   :   assert (rdbk == 32'h0000001e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	267   :   assert (rdbk == 32'h000000da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	268   :   assert (rdbk == 32'h000000f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	269   :   assert (rdbk == 32'h00000058) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	270   :   assert (rdbk == 32'hffffff0e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	271   :   assert (rdbk == 32'h000000c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	272   :   assert (rdbk == 32'hfffffff2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	273   :   assert (rdbk == 32'hffffff29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	274   :   assert (rdbk == 32'h000000a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	275   :   assert (rdbk == 32'hffffff77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	276   :   assert (rdbk == 32'hffffffc1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	277   :   assert (rdbk == 32'h0000001b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	278   :   assert (rdbk == 32'h0000003d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	279   :   assert (rdbk == 32'h00000052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	280   :   assert (rdbk == 32'h0000009e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	281   :   assert (rdbk == 32'hffffff95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	282   :   assert (rdbk == 32'h0000004d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	283   :   assert (rdbk == 32'hfffffeb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	284   :   assert (rdbk == 32'h00000053) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	285   :   assert (rdbk == 32'hfffffee0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	286   :   assert (rdbk == 32'hffffffc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	287   :   assert (rdbk == 32'hffffffcc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	288   :   assert (rdbk == 32'hffffff29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	289   :   assert (rdbk == 32'h0000006e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	290   :   assert (rdbk == 32'h00000024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	291   :   assert (rdbk == 32'h000000f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	292   :   assert (rdbk == 32'hffffffe1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	293   :   assert (rdbk == 32'hffffff2a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	294   :   assert (rdbk == 32'h0000008f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	295   :   assert (rdbk == 32'h0000002d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	296   :   assert (rdbk == 32'h00000056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	297   :   assert (rdbk == 32'hffffff2f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	298   :   assert (rdbk == 32'hffffff35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	299   :   assert (rdbk == 32'h00000025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	300   :   assert (rdbk == 32'hffffff4c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	301   :   assert (rdbk == 32'h00000026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	302   :   assert (rdbk == 32'hffffff26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	303   :   assert (rdbk == 32'h000000c4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	304   :   assert (rdbk == 32'hffffff5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	305   :   assert (rdbk == 32'h000000ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	306   :   assert (rdbk == 32'hffffffc2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	307   :   assert (rdbk == 32'hffffff6a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	308   :   assert (rdbk == 32'hffffffd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	309   :   assert (rdbk == 32'h00000081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	310   :   assert (rdbk == 32'hffffff6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	311   :   assert (rdbk == 32'hffffff64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	312   :   assert (rdbk == 32'hffffff7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	313   :   assert (rdbk == 32'hffffffc1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	314   :   assert (rdbk == 32'hffffff93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	315   :   assert (rdbk == 32'hffffffaf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	316   :   assert (rdbk == 32'hffffffa6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	317   :   assert (rdbk == 32'hffffff9d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	318   :   assert (rdbk == 32'h000000a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	319   :   assert (rdbk == 32'hffffff7b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	320   :   assert (rdbk == 32'h0000008f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	321   :   assert (rdbk == 32'hfffffff7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	322   :   assert (rdbk == 32'hffffffc7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	323   :   assert (rdbk == 32'h0000001f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	324   :   assert (rdbk == 32'hfffffff8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	325   :   assert (rdbk == 32'h00000061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	326   :   assert (rdbk == 32'hffffff0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	327   :   assert (rdbk == 32'hffffffb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	328   :   assert (rdbk == 32'h000000d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	329   :   assert (rdbk == 32'h00000099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	330   :   assert (rdbk == 32'h00000046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	331   :   assert (rdbk == 32'h0000000d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	332   :   assert (rdbk == 32'h00000088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	333   :   assert (rdbk == 32'h000000bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	334   :   assert (rdbk == 32'h00000007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	335   :   assert (rdbk == 32'hfffffed5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	336   :   assert (rdbk == 32'h0000001b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	337   :   assert (rdbk == 32'h0000004b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	338   :   assert (rdbk == 32'h00000086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	339   :   assert (rdbk == 32'hffffff59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	340   :   assert (rdbk == 32'h0000003a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	341   :   assert (rdbk == 32'h00000015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	342   :   assert (rdbk == 32'hfffffff4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	343   :   assert (rdbk == 32'h0000004b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	344   :   assert (rdbk == 32'hffffff83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	345   :   assert (rdbk == 32'hffffffc6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	346   :   assert (rdbk == 32'h00000098) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	347   :   assert (rdbk == 32'hffffffd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	348   :   assert (rdbk == 32'hfffffffc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	349   :   assert (rdbk == 32'h00000018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	350   :   assert (rdbk == 32'h00000150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	351   :   assert (rdbk == 32'hffffffae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	352   :   assert (rdbk == 32'hffffff38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	353   :   assert (rdbk == 32'h0000000f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	354   :   assert (rdbk == 32'hffffff33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	355   :   assert (rdbk == 32'h000000f8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	356   :   assert (rdbk == 32'h000000bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	357   :   assert (rdbk == 32'hffffff76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	358   :   assert (rdbk == 32'hffffffee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	359   :   assert (rdbk == 32'hfffffeca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	360   :   assert (rdbk == 32'h00000067) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	361   :   assert (rdbk == 32'hffffff5c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	362   :   assert (rdbk == 32'h0000002c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	363   :   assert (rdbk == 32'h00000050) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	364   :   assert (rdbk == 32'hffffffdb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	365   :   assert (rdbk == 32'h00000043) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	366   :   assert (rdbk == 32'hffffff9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	367   :   assert (rdbk == 32'hffffffce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	368   :   assert (rdbk == 32'h0000003b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	369   :   assert (rdbk == 32'hffffff5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	370   :   assert (rdbk == 32'hffffffb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	371   :   assert (rdbk == 32'h000000a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	372   :   assert (rdbk == 32'hffffff24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	373   :   assert (rdbk == 32'hffffff39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	374   :   assert (rdbk == 32'h00000122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	375   :   assert (rdbk == 32'h00000083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	376   :   assert (rdbk == 32'hffffffaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	377   :   assert (rdbk == 32'hfffffea2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	378   :   assert (rdbk == 32'hffffff62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	379   :   assert (rdbk == 32'hfffffff4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	380   :   assert (rdbk == 32'h00000018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	381   :   assert (rdbk == 32'h000000aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	382   :   assert (rdbk == 32'hffffffb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	383   :   assert (rdbk == 32'h0000012b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	384   :   assert (rdbk == 32'h00000006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	385   :   assert (rdbk == 32'h00000017) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	386   :   assert (rdbk == 32'hffffffdf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	387   :   assert (rdbk == 32'hffffff71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	388   :   assert (rdbk == 32'h00000038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	389   :   assert (rdbk == 32'h00000046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	390   :   assert (rdbk == 32'h000000c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	391   :   assert (rdbk == 32'hffffffc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	392   :   assert (rdbk == 32'hffffffee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	393   :   assert (rdbk == 32'hfffffffd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	394   :   assert (rdbk == 32'hffffffd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	395   :   assert (rdbk == 32'h00000091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	396   :   assert (rdbk == 32'h0000000a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	397   :   assert (rdbk == 32'hffffffae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	398   :   assert (rdbk == 32'h00000224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	399   :   assert (rdbk == 32'hffffffc2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	400   :   assert (rdbk == 32'h00000163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	401   :   assert (rdbk == 32'h00000091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	402   :   assert (rdbk == 32'hfffffff5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	403   :   assert (rdbk == 32'hffffff86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	404   :   assert (rdbk == 32'h000000b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	405   :   assert (rdbk == 32'h000000cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	406   :   assert (rdbk == 32'h00000026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	407   :   assert (rdbk == 32'h00000073) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	408   :   assert (rdbk == 32'hffffff35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	409   :   assert (rdbk == 32'h00000091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	410   :   assert (rdbk == 32'hfffffee9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	411   :   assert (rdbk == 32'hffffff09) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	412   :   assert (rdbk == 32'hffffff9e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	413   :   assert (rdbk == 32'h00000066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	414   :   assert (rdbk == 32'h0000001c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	415   :   assert (rdbk == 32'h00000058) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	416   :   assert (rdbk == 32'h0000003b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	417   :   assert (rdbk == 32'h00000190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	418   :   assert (rdbk == 32'hffffffa3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	419   :   assert (rdbk == 32'h00000067) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	420   :   assert (rdbk == 32'h00000098) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	421   :   assert (rdbk == 32'hffffff83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	422   :   assert (rdbk == 32'hffffff75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	423   :   assert (rdbk == 32'h00000060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	424   :   assert (rdbk == 32'h00000071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	425   :   assert (rdbk == 32'hffffffb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	426   :   assert (rdbk == 32'h0000002a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	427   :   assert (rdbk == 32'h00000050) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	428   :   assert (rdbk == 32'hfffffffc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	429   :   assert (rdbk == 32'hffffffb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	430   :   assert (rdbk == 32'h00000035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	431   :   assert (rdbk == 32'hfffffedd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	432   :   assert (rdbk == 32'h00000053) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	433   :   assert (rdbk == 32'h000000a4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	434   :   assert (rdbk == 32'hfffffee0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	435   :   assert (rdbk == 32'hffffffc1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	436   :   assert (rdbk == 32'h000000b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	437   :   assert (rdbk == 32'hffffffbb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	438   :   assert (rdbk == 32'hffffff5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	439   :   assert (rdbk == 32'h00000026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	440   :   assert (rdbk == 32'h00000089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	441   :   assert (rdbk == 32'hfffffee8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	442   :   assert (rdbk == 32'h00000008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	443   :   assert (rdbk == 32'h0000006b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	444   :   assert (rdbk == 32'h000000e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	445   :   assert (rdbk == 32'hffffffe7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	446   :   assert (rdbk == 32'h0000001c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	447   :   assert (rdbk == 32'h000000fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	448   :   assert (rdbk == 32'h000000ae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	449   :   assert (rdbk == 32'h0000003d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	450   :   assert (rdbk == 32'h000000be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	451   :   assert (rdbk == 32'h000000d9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	452   :   assert (rdbk == 32'h000000c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	453   :   assert (rdbk == 32'h0000001e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	454   :   assert (rdbk == 32'hffffff82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	455   :   assert (rdbk == 32'hffffff2f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	456   :   assert (rdbk == 32'hffffffda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	457   :   assert (rdbk == 32'hffffff72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	458   :   assert (rdbk == 32'h0000009e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	459   :   assert (rdbk == 32'h0000013d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	460   :   assert (rdbk == 32'hfffffff9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	461   :   assert (rdbk == 32'hffffffde) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	462   :   assert (rdbk == 32'h00000021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	463   :   assert (rdbk == 32'h00000063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	464   :   assert (rdbk == 32'h00000051) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	465   :   assert (rdbk == 32'h0000001c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	466   :   assert (rdbk == 32'hffffff78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	467   :   assert (rdbk == 32'hffffff77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	468   :   assert (rdbk == 32'hffffff2b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	469   :   assert (rdbk == 32'h00000027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	470   :   assert (rdbk == 32'h00000013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	471   :   assert (rdbk == 32'h000001c4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	472   :   assert (rdbk == 32'h0000003c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	473   :   assert (rdbk == 32'hffffffeb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	474   :   assert (rdbk == 32'hffffff31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	475   :   assert (rdbk == 32'hffffffa2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	476   :   assert (rdbk == 32'hfffffe5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	477   :   assert (rdbk == 32'h00000013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	478   :   assert (rdbk == 32'hffffff13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	479   :   assert (rdbk == 32'h00000015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	480   :   assert (rdbk == 32'hffffff11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	481   :   assert (rdbk == 32'h000000b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	482   :   assert (rdbk == 32'hffffff79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	483   :   assert (rdbk == 32'h000000a9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	484   :   assert (rdbk == 32'h0000002f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	485   :   assert (rdbk == 32'h00000053) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	486   :   assert (rdbk == 32'h00000110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	487   :   assert (rdbk == 32'hfffffe64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	488   :   assert (rdbk == 32'h00000056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	489   :   assert (rdbk == 32'h00000047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	490   :   assert (rdbk == 32'hfffffebb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	491   :   assert (rdbk == 32'h000000a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	492   :   assert (rdbk == 32'hfffffe8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	493   :   assert (rdbk == 32'h00000038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	494   :   assert (rdbk == 32'hffffff90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	495   :   assert (rdbk == 32'h00000041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	496   :   assert (rdbk == 32'h000000b2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	497   :   assert (rdbk == 32'hffffffe0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	498   :   assert (rdbk == 32'hffffffd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	499   :   assert (rdbk == 32'h00000145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	500   :   assert (rdbk == 32'h00000064) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	501   :   assert (rdbk == 32'hfffffea2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	502   :   assert (rdbk == 32'h00000177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	503   :   assert (rdbk == 32'hffffffa3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	504   :   assert (rdbk == 32'h00000061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	505   :   assert (rdbk == 32'h000000c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	506   :   assert (rdbk == 32'hfffffe66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	507   :   assert (rdbk == 32'hffffff62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	508   :   assert (rdbk == 32'h000000ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	509   :   assert (rdbk == 32'hffffffe6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	510   :   assert (rdbk == 32'hfffffecb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	511   :   assert (rdbk == 32'hffffff90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	512   :   assert (rdbk == 32'h000000b2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	513   :   assert (rdbk == 32'h0000000b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	514   :   assert (rdbk == 32'hffffff99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	515   :   assert (rdbk == 32'hfffffdd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	516   :   assert (rdbk == 32'h0000004f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	517   :   assert (rdbk == 32'h00000076) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	518   :   assert (rdbk == 32'h000000ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	519   :   assert (rdbk == 32'h000000dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	520   :   assert (rdbk == 32'h00000078) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	521   :   assert (rdbk == 32'hffffff66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	522   :   assert (rdbk == 32'h00000002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	523   :   assert (rdbk == 32'h00000007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	524   :   assert (rdbk == 32'hffffff05) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	525   :   assert (rdbk == 32'hffffffa3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	526   :   assert (rdbk == 32'hfffffff7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	527   :   assert (rdbk == 32'h00000010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	528   :   assert (rdbk == 32'h0000004a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	529   :   assert (rdbk == 32'h00000072) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	530   :   assert (rdbk == 32'hffffffda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	531   :   assert (rdbk == 32'h000000a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	532   :   assert (rdbk == 32'h00000073) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	533   :   assert (rdbk == 32'h000000ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	534   :   assert (rdbk == 32'hfffffff2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	535   :   assert (rdbk == 32'hffffff66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	536   :   assert (rdbk == 32'h00000075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	537   :   assert (rdbk == 32'hffffff9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	538   :   assert (rdbk == 32'hffffff69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	539   :   assert (rdbk == 32'hffffff3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	540   :   assert (rdbk == 32'hffffff60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	541   :   assert (rdbk == 32'h0000003b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	542   :   assert (rdbk == 32'h0000006e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	543   :   assert (rdbk == 32'h000001d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	544   :   assert (rdbk == 32'h00000121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	545   :   assert (rdbk == 32'hffffff77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	546   :   assert (rdbk == 32'hffffff66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	547   :   assert (rdbk == 32'hffffff40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	548   :   assert (rdbk == 32'hfffffef3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	549   :   assert (rdbk == 32'h00000108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	550   :   assert (rdbk == 32'h0000001b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	551   :   assert (rdbk == 32'h000000d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	552   :   assert (rdbk == 32'h0000004c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	553   :   assert (rdbk == 32'h00000075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	554   :   assert (rdbk == 32'hffffffca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	555   :   assert (rdbk == 32'h000000d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	556   :   assert (rdbk == 32'h000000fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	557   :   assert (rdbk == 32'h000000b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	558   :   assert (rdbk == 32'h000000dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	559   :   assert (rdbk == 32'hffffff03) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	560   :   assert (rdbk == 32'h00000041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	561   :   assert (rdbk == 32'hffffff08) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	562   :   assert (rdbk == 32'hffffff41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	563   :   assert (rdbk == 32'h0000000b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	564   :   assert (rdbk == 32'h00000084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	565   :   assert (rdbk == 32'hffffff42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	566   :   assert (rdbk == 32'hffffffcc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	567   :   assert (rdbk == 32'hffffffad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	568   :   assert (rdbk == 32'h00000063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	569   :   assert (rdbk == 32'hffffff89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	570   :   assert (rdbk == 32'h0000009b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	571   :   assert (rdbk == 32'h0000008b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	572   :   assert (rdbk == 32'hfffffff2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	573   :   assert (rdbk == 32'hffffffc8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	574   :   assert (rdbk == 32'hffffffdd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	575   :   assert (rdbk == 32'hffffff61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	576   :   assert (rdbk == 32'hffffffab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	577   :   assert (rdbk == 32'h000000b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	578   :   assert (rdbk == 32'h00000026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	579   :   assert (rdbk == 32'h000000dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	580   :   assert (rdbk == 32'hffffff44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	581   :   assert (rdbk == 32'hffffff91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	582   :   assert (rdbk == 32'h000000bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	583   :   assert (rdbk == 32'h0000001e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	584   :   assert (rdbk == 32'hffffffe3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	585   :   assert (rdbk == 32'h00000018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	586   :   assert (rdbk == 32'hffffff37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	587   :   assert (rdbk == 32'h0000017d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	588   :   assert (rdbk == 32'hffffff8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	589   :   assert (rdbk == 32'hffffff38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	590   :   assert (rdbk == 32'h00000012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	591   :   assert (rdbk == 32'h00000035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	592   :   assert (rdbk == 32'h00000035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	593   :   assert (rdbk == 32'h000000cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	594   :   assert (rdbk == 32'hfffffeee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	595   :   assert (rdbk == 32'h00000059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	596   :   assert (rdbk == 32'hffffff96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	597   :   assert (rdbk == 32'h00000173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	598   :   assert (rdbk == 32'hffffffc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	599   :   assert (rdbk == 32'h000000b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	600   :   assert (rdbk == 32'h00000011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	601   :   assert (rdbk == 32'h000000bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	602   :   assert (rdbk == 32'hfffffe3b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	603   :   assert (rdbk == 32'hffffff41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	604   :   assert (rdbk == 32'hffffff5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	605   :   assert (rdbk == 32'h00000013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	606   :   assert (rdbk == 32'h0000015b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	607   :   assert (rdbk == 32'hffffff9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	608   :   assert (rdbk == 32'h0000002d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	609   :   assert (rdbk == 32'hffffffbe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	610   :   assert (rdbk == 32'h00000093) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	611   :   assert (rdbk == 32'hfffffed5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	612   :   assert (rdbk == 32'hffffffbd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	613   :   assert (rdbk == 32'hffffff29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	614   :   assert (rdbk == 32'hffffffb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	615   :   assert (rdbk == 32'h00000189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	616   :   assert (rdbk == 32'hfffffeac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	617   :   assert (rdbk == 32'h00000069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	618   :   assert (rdbk == 32'h0000007e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	619   :   assert (rdbk == 32'hffffffc6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	620   :   assert (rdbk == 32'h00000084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	621   :   assert (rdbk == 32'hffffff31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	622   :   assert (rdbk == 32'hffffff5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	623   :   assert (rdbk == 32'hffffff88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	624   :   assert (rdbk == 32'hfffffdff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	625   :   assert (rdbk == 32'hffffff23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	626   :   assert (rdbk == 32'h0000000c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	627   :   assert (rdbk == 32'h000000c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	628   :   assert (rdbk == 32'h0000007d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	629   :   assert (rdbk == 32'hffffff94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	630   :   assert (rdbk == 32'hffffff90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	631   :   assert (rdbk == 32'h0000002b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	632   :   assert (rdbk == 32'hffffffdd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	633   :   assert (rdbk == 32'hffffff4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	634   :   assert (rdbk == 32'hffffffe5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	635   :   assert (rdbk == 32'h0000009d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	636   :   assert (rdbk == 32'hffffffed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	637   :   assert (rdbk == 32'h00000067) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	638   :   assert (rdbk == 32'h00000004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	639   :   assert (rdbk == 32'hffffff9c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	640   :   assert (rdbk == 32'hffffffab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	641   :   assert (rdbk == 32'hffffff4c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	642   :   assert (rdbk == 32'h000000af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	643   :   assert (rdbk == 32'h00000101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	644   :   assert (rdbk == 32'h00000027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	645   :   assert (rdbk == 32'h000000d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	646   :   assert (rdbk == 32'hffffff6a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	647   :   assert (rdbk == 32'h00000001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	648   :   assert (rdbk == 32'h000000f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	649   :   assert (rdbk == 32'h00000022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	650   :   assert (rdbk == 32'hffffff5c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	651   :   assert (rdbk == 32'h00000028) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	652   :   assert (rdbk == 32'h000000d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	653   :   assert (rdbk == 32'h00000037) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	654   :   assert (rdbk == 32'h00000056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	655   :   assert (rdbk == 32'hfffffed0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	656   :   assert (rdbk == 32'h00000085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	657   :   assert (rdbk == 32'hffffff94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	658   :   assert (rdbk == 32'h000000e2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	659   :   assert (rdbk == 32'hffffff8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	660   :   assert (rdbk == 32'hffffff9c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	661   :   assert (rdbk == 32'h00000056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	662   :   assert (rdbk == 32'hffffff47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	663   :   assert (rdbk == 32'hffffff8c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	664   :   assert (rdbk == 32'hffffff28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	665   :   assert (rdbk == 32'hffffffa2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	666   :   assert (rdbk == 32'h00000111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	667   :   assert (rdbk == 32'hffffff9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	668   :   assert (rdbk == 32'hffffffca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	669   :   assert (rdbk == 32'h000000f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	670   :   assert (rdbk == 32'h000001b1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	671   :   assert (rdbk == 32'hffffffcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	672   :   assert (rdbk == 32'h000000fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	673   :   assert (rdbk == 32'h000000fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	674   :   assert (rdbk == 32'h0000001d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	675   :   assert (rdbk == 32'hffffff94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	676   :   assert (rdbk == 32'hffffff4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	677   :   assert (rdbk == 32'h00000074) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	678   :   assert (rdbk == 32'hffffffd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	679   :   assert (rdbk == 32'h000000ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	680   :   assert (rdbk == 32'h000000a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	681   :   assert (rdbk == 32'hffffff9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	682   :   assert (rdbk == 32'hffffffe3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	683   :   assert (rdbk == 32'hfffffefc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	684   :   assert (rdbk == 32'h0000006d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	685   :   assert (rdbk == 32'h0000001c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	686   :   assert (rdbk == 32'h00000082) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	687   :   assert (rdbk == 32'hffffff76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	688   :   assert (rdbk == 32'hffffff96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	689   :   assert (rdbk == 32'h00000073) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	690   :   assert (rdbk == 32'hffffff15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	691   :   assert (rdbk == 32'h00000004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	692   :   assert (rdbk == 32'h00000002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	693   :   assert (rdbk == 32'hffffffb1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	694   :   assert (rdbk == 32'hffffff35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	695   :   assert (rdbk == 32'h00000011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	696   :   assert (rdbk == 32'h0000006b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	697   :   assert (rdbk == 32'hffffffe8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	698   :   assert (rdbk == 32'hffffff2b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	699   :   assert (rdbk == 32'h0000007c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	700   :   assert (rdbk == 32'hfffffffe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	701   :   assert (rdbk == 32'hffffffd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	702   :   assert (rdbk == 32'hffffffa7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	703   :   assert (rdbk == 32'h00000079) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	704   :   assert (rdbk == 32'h0000005e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	705   :   assert (rdbk == 32'hfffffe9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	706   :   assert (rdbk == 32'h00000072) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	707   :   assert (rdbk == 32'hffffff77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	708   :   assert (rdbk == 32'hffffff07) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	709   :   assert (rdbk == 32'h00000094) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	710   :   assert (rdbk == 32'hfffffff9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	711   :   assert (rdbk == 32'h0000009c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	712   :   assert (rdbk == 32'hffffff60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	713   :   assert (rdbk == 32'hffffff9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	714   :   assert (rdbk == 32'hffffffb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	715   :   assert (rdbk == 32'hfffffef1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	716   :   assert (rdbk == 32'hffffffbb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	717   :   assert (rdbk == 32'h00000035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	718   :   assert (rdbk == 32'h0000002e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	719   :   assert (rdbk == 32'hffffffcd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	720   :   assert (rdbk == 32'h00000066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	721   :   assert (rdbk == 32'hfffffff2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	722   :   assert (rdbk == 32'hffffff22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	723   :   assert (rdbk == 32'h00000014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	724   :   assert (rdbk == 32'hfffffe91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	725   :   assert (rdbk == 32'h0000007d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	726   :   assert (rdbk == 32'h00000104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	727   :   assert (rdbk == 32'hffffffff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	728   :   assert (rdbk == 32'h000000a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	729   :   assert (rdbk == 32'h00000021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	730   :   assert (rdbk == 32'h0000011e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	731   :   assert (rdbk == 32'h000000c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	732   :   assert (rdbk == 32'h00000023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	733   :   assert (rdbk == 32'h0000007c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	734   :   assert (rdbk == 32'hffffff37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	735   :   assert (rdbk == 32'h00000072) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	736   :   assert (rdbk == 32'hffffffba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	737   :   assert (rdbk == 32'h00000030) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	738   :   assert (rdbk == 32'hffffffbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	739   :   assert (rdbk == 32'h00000057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	740   :   assert (rdbk == 32'h000000ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	741   :   assert (rdbk == 32'hffffffa3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	742   :   assert (rdbk == 32'h0000002f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	743   :   assert (rdbk == 32'hffffff41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	744   :   assert (rdbk == 32'h0000001d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	745   :   assert (rdbk == 32'h00000099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	746   :   assert (rdbk == 32'h000000ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	747   :   assert (rdbk == 32'h00000135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	748   :   assert (rdbk == 32'h0000012c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	749   :   assert (rdbk == 32'hfffffff8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	750   :   assert (rdbk == 32'hffffffc4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	751   :   assert (rdbk == 32'hffffff79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	752   :   assert (rdbk == 32'hffffff70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	753   :   assert (rdbk == 32'h0000010f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	754   :   assert (rdbk == 32'h0000000d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	755   :   assert (rdbk == 32'hfffffff1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	756   :   assert (rdbk == 32'h000000f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	757   :   assert (rdbk == 32'hffffffda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	758   :   assert (rdbk == 32'hffffff86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	759   :   assert (rdbk == 32'h0000013d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	760   :   assert (rdbk == 32'h0000000f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	761   :   assert (rdbk == 32'hfffffec4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	762   :   assert (rdbk == 32'hfffffe77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	763   :   assert (rdbk == 32'h00000078) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	764   :   assert (rdbk == 32'hffffffc7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	765   :   assert (rdbk == 32'h0000000c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	766   :   assert (rdbk == 32'hffffffcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	767   :   assert (rdbk == 32'hffffff54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	768   :   assert (rdbk == 32'hffffff48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	769   :   assert (rdbk == 32'h000000af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	770   :   assert (rdbk == 32'hffffff5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	771   :   assert (rdbk == 32'hffffff39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	772   :   assert (rdbk == 32'hffffff6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	773   :   assert (rdbk == 32'h00000050) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	774   :   assert (rdbk == 32'hfffffff5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	775   :   assert (rdbk == 32'hfffffee0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	776   :   assert (rdbk == 32'hfffffefe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	777   :   assert (rdbk == 32'hffffffd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	778   :   assert (rdbk == 32'h0000004e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	779   :   assert (rdbk == 32'hffffffdd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	780   :   assert (rdbk == 32'hffffff1e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	781   :   assert (rdbk == 32'hffffff97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	782   :   assert (rdbk == 32'h00000047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	783   :   assert (rdbk == 32'h00000123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	784   :   assert (rdbk == 32'h0000003b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	785   :   assert (rdbk == 32'hffffff3f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	786   :   assert (rdbk == 32'hffffff63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	787   :   assert (rdbk == 32'hffffffca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	788   :   assert (rdbk == 32'hffffff30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	789   :   assert (rdbk == 32'h0000004a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	790   :   assert (rdbk == 32'h00000086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	791   :   assert (rdbk == 32'hffffff64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	792   :   assert (rdbk == 32'h00000078) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	793   :   assert (rdbk == 32'h000000a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	794   :   assert (rdbk == 32'hffffff26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	795   :   assert (rdbk == 32'hffffff3e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	796   :   assert (rdbk == 32'h00000065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	797   :   assert (rdbk == 32'h0000001f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	798   :   assert (rdbk == 32'hffffffdd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	799   :   assert (rdbk == 32'hffffff72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	800   :   assert (rdbk == 32'h0000009c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	801   :   assert (rdbk == 32'hfffffece) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	802   :   assert (rdbk == 32'hffffffa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	803   :   assert (rdbk == 32'h00000101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	804   :   assert (rdbk == 32'hffffff23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	805   :   assert (rdbk == 32'h000000af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	806   :   assert (rdbk == 32'hffffffe5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	807   :   assert (rdbk == 32'hffffff15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	808   :   assert (rdbk == 32'hfffffff1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	809   :   assert (rdbk == 32'h0000011e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	810   :   assert (rdbk == 32'h0000001b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	811   :   assert (rdbk == 32'h000000b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	812   :   assert (rdbk == 32'hffffff3d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	813   :   assert (rdbk == 32'h0000002e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	814   :   assert (rdbk == 32'h000000b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	815   :   assert (rdbk == 32'h000000f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	816   :   assert (rdbk == 32'hfffffffa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	817   :   assert (rdbk == 32'hffffff9c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	818   :   assert (rdbk == 32'h00000026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	819   :   assert (rdbk == 32'h00000059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	820   :   assert (rdbk == 32'h000000ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	821   :   assert (rdbk == 32'h00000106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	822   :   assert (rdbk == 32'h00000149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	823   :   assert (rdbk == 32'hffffff67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	824   :   assert (rdbk == 32'hffffff11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	825   :   assert (rdbk == 32'h00000012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	826   :   assert (rdbk == 32'h00000077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	827   :   assert (rdbk == 32'h000000fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	828   :   assert (rdbk == 32'h00000011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	829   :   assert (rdbk == 32'h0000006e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	830   :   assert (rdbk == 32'h00000062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	831   :   assert (rdbk == 32'hffffff89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	832   :   assert (rdbk == 32'h00000127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	833   :   assert (rdbk == 32'h0000000e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	834   :   assert (rdbk == 32'h00000020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	835   :   assert (rdbk == 32'h00000207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	836   :   assert (rdbk == 32'h00000081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	837   :   assert (rdbk == 32'h0000005a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	838   :   assert (rdbk == 32'h0000004b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	839   :   assert (rdbk == 32'h000000c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	840   :   assert (rdbk == 32'hfffffedf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	841   :   assert (rdbk == 32'hfffffef0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	842   :   assert (rdbk == 32'h00000035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	843   :   assert (rdbk == 32'h0000006d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	844   :   assert (rdbk == 32'hffffff95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	845   :   assert (rdbk == 32'h0000017d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	846   :   assert (rdbk == 32'h00000011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	847   :   assert (rdbk == 32'h000000dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	848   :   assert (rdbk == 32'hfffffff2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	849   :   assert (rdbk == 32'h00000008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	850   :   assert (rdbk == 32'hffffff6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	851   :   assert (rdbk == 32'hffffff73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	852   :   assert (rdbk == 32'h0000004d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	853   :   assert (rdbk == 32'h00000021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	854   :   assert (rdbk == 32'h00000094) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	855   :   assert (rdbk == 32'hfffffebb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	856   :   assert (rdbk == 32'h000000b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	857   :   assert (rdbk == 32'h00000005) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	858   :   assert (rdbk == 32'hffffffad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	859   :   assert (rdbk == 32'h0000000a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	860   :   assert (rdbk == 32'h000000be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	861   :   assert (rdbk == 32'h0000009b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	862   :   assert (rdbk == 32'h00000164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	863   :   assert (rdbk == 32'h00000056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	864   :   assert (rdbk == 32'hffffffe6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	865   :   assert (rdbk == 32'hffffff18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	866   :   assert (rdbk == 32'h00000051) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	867   :   assert (rdbk == 32'hffffff6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	868   :   assert (rdbk == 32'h000000c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	869   :   assert (rdbk == 32'h0000001c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	870   :   assert (rdbk == 32'hfffffe82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	871   :   assert (rdbk == 32'hffffffa2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	872   :   assert (rdbk == 32'hffffff36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	873   :   assert (rdbk == 32'h000000c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	874   :   assert (rdbk == 32'h0000009b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	875   :   assert (rdbk == 32'h00000184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	876   :   assert (rdbk == 32'hfffffe21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	877   :   assert (rdbk == 32'hffffff4e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	878   :   assert (rdbk == 32'h000000d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	879   :   assert (rdbk == 32'hffffffcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	880   :   assert (rdbk == 32'hffffffba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	881   :   assert (rdbk == 32'hffffffca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	882   :   assert (rdbk == 32'h00000085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	883   :   assert (rdbk == 32'h0000006e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	884   :   assert (rdbk == 32'h000000e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	885   :   assert (rdbk == 32'h000000da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	886   :   assert (rdbk == 32'hffffffdb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	887   :   assert (rdbk == 32'hfffffeda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	888   :   assert (rdbk == 32'h00000062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	889   :   assert (rdbk == 32'hffffffac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	890   :   assert (rdbk == 32'h00000049) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	891   :   assert (rdbk == 32'h00000098) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	892   :   assert (rdbk == 32'hffffffc7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	893   :   assert (rdbk == 32'hffffffba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	894   :   assert (rdbk == 32'hffffff91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	895   :   assert (rdbk == 32'hffffff8d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	896   :   assert (rdbk == 32'hffffff6a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	897   :   assert (rdbk == 32'h000000c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	898   :   assert (rdbk == 32'h00000037) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	899   :   assert (rdbk == 32'h00000094) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	900   :   assert (rdbk == 32'h000000ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	901   :   assert (rdbk == 32'h000000b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	902   :   assert (rdbk == 32'h00000014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	903   :   assert (rdbk == 32'hfffffe9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	904   :   assert (rdbk == 32'h000000ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	905   :   assert (rdbk == 32'hffffff41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	906   :   assert (rdbk == 32'h0000001e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	907   :   assert (rdbk == 32'hffffffc0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	908   :   assert (rdbk == 32'h00000089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	909   :   assert (rdbk == 32'h00000000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	910   :   assert (rdbk == 32'hffffffa6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	911   :   assert (rdbk == 32'h0000000a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	912   :   assert (rdbk == 32'hffffffe5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	913   :   assert (rdbk == 32'h00000014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	914   :   assert (rdbk == 32'hffffffb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	915   :   assert (rdbk == 32'h00000104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	916   :   assert (rdbk == 32'hffffffb7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	917   :   assert (rdbk == 32'h0000008e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	918   :   assert (rdbk == 32'hffffffde) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	919   :   assert (rdbk == 32'hffffff4e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	920   :   assert (rdbk == 32'h00000006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	921   :   assert (rdbk == 32'hffffff8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	922   :   assert (rdbk == 32'hffffff02) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	923   :   assert (rdbk == 32'hfffffe9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	924   :   assert (rdbk == 32'h00000000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	925   :   assert (rdbk == 32'hffffff84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	926   :   assert (rdbk == 32'h0000001d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	927   :   assert (rdbk == 32'h0000005a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	928   :   assert (rdbk == 32'h0000009c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	929   :   assert (rdbk == 32'h00000120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	930   :   assert (rdbk == 32'hfffffff2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	931   :   assert (rdbk == 32'hfffffffd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	932   :   assert (rdbk == 32'hffffffec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	933   :   assert (rdbk == 32'h0000008e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	934   :   assert (rdbk == 32'hfffffff8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	935   :   assert (rdbk == 32'hffffff46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	936   :   assert (rdbk == 32'hffffff85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	937   :   assert (rdbk == 32'hffffff95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	938   :   assert (rdbk == 32'h0000010d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	939   :   assert (rdbk == 32'h0000005b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	940   :   assert (rdbk == 32'h0000019d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	941   :   assert (rdbk == 32'h00000085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	942   :   assert (rdbk == 32'hfffffffb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	943   :   assert (rdbk == 32'h0000002e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	944   :   assert (rdbk == 32'hfffffefb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	945   :   assert (rdbk == 32'hffffffd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	946   :   assert (rdbk == 32'h00000085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	947   :   assert (rdbk == 32'hffffff91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	948   :   assert (rdbk == 32'hffffff92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	949   :   assert (rdbk == 32'h00000013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	950   :   assert (rdbk == 32'h0000003b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	951   :   assert (rdbk == 32'h0000008a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	952   :   assert (rdbk == 32'h00000002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	953   :   assert (rdbk == 32'h00000036) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	954   :   assert (rdbk == 32'hfffffe1a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	955   :   assert (rdbk == 32'h0000006a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	956   :   assert (rdbk == 32'hffffffd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	957   :   assert (rdbk == 32'hffffff34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	958   :   assert (rdbk == 32'h0000010e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	959   :   assert (rdbk == 32'h00000086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	960   :   assert (rdbk == 32'h00000118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	961   :   assert (rdbk == 32'hffffffb6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	962   :   assert (rdbk == 32'hfffffe64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	963   :   assert (rdbk == 32'hfffffe86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	964   :   assert (rdbk == 32'hfffffeaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	965   :   assert (rdbk == 32'hffffff7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	966   :   assert (rdbk == 32'h0000009a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	967   :   assert (rdbk == 32'hffffff52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	968   :   assert (rdbk == 32'h00000019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	969   :   assert (rdbk == 32'hffffff9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	970   :   assert (rdbk == 32'h000000d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	971   :   assert (rdbk == 32'hffffff28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	972   :   assert (rdbk == 32'h000001a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	973   :   assert (rdbk == 32'h0000019e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	974   :   assert (rdbk == 32'h000000a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	975   :   assert (rdbk == 32'h00000015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	976   :   assert (rdbk == 32'h00000104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	977   :   assert (rdbk == 32'h0000006e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	978   :   assert (rdbk == 32'h000000be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	979   :   assert (rdbk == 32'hffffff82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	980   :   assert (rdbk == 32'hfffffff5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	981   :   assert (rdbk == 32'hffffff9e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	982   :   assert (rdbk == 32'hffffffa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	983   :   assert (rdbk == 32'h000000a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	984   :   assert (rdbk == 32'hffffff87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	985   :   assert (rdbk == 32'hffffff2d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	986   :   assert (rdbk == 32'hffffffd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	987   :   assert (rdbk == 32'hfffffff3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	988   :   assert (rdbk == 32'hfffffe9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	989   :   assert (rdbk == 32'h00000048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	990   :   assert (rdbk == 32'hffffff73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	991   :   assert (rdbk == 32'hffffffcd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	992   :   assert (rdbk == 32'h00000093) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	993   :   assert (rdbk == 32'hfffffeda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	994   :   assert (rdbk == 32'h0000006b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	995   :   assert (rdbk == 32'h000000f8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	996   :   assert (rdbk == 32'hffffffbc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	997   :   assert (rdbk == 32'hffffff31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	998   :   assert (rdbk == 32'h00000090) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	999   :   assert (rdbk == 32'hffffff68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1000   :   assert (rdbk == 32'hffffff66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1001   :   assert (rdbk == 32'hffffff36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1002   :   assert (rdbk == 32'hffffffc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1003   :   assert (rdbk == 32'h0000008f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1004   :   assert (rdbk == 32'h00000091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1005   :   assert (rdbk == 32'h00000076) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1006   :   assert (rdbk == 32'h0000000f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1007   :   assert (rdbk == 32'hfffffff4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1008   :   assert (rdbk == 32'hffffff33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1009   :   assert (rdbk == 32'hffffff8e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1010   :   assert (rdbk == 32'h00000003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1011   :   assert (rdbk == 32'hffffffdb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1012   :   assert (rdbk == 32'hffffff9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1013   :   assert (rdbk == 32'hffffffc0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1014   :   assert (rdbk == 32'hffffff78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1015   :   assert (rdbk == 32'h00000018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1016   :   assert (rdbk == 32'hffffffa5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1017   :   assert (rdbk == 32'h00000034) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1018   :   assert (rdbk == 32'hfffffff3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1019   :   assert (rdbk == 32'hfffffe69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1020   :   assert (rdbk == 32'h000000d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1021   :   assert (rdbk == 32'h00000010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1022   :   assert (rdbk == 32'hffffffe2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1023   :   assert (rdbk == 32'h0000003f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
endcase
end

