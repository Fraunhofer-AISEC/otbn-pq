// Copyright Copyright Fraunhofer Institute for Applied and Integrated Security (AISEC).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

$fwrite(f,"----------------------------------------------------------------\n");   
$fwrite(f,"-- PQ-INVNTT-Indirect (Falcon-1024)\n");
$fwrite(f,"----------------------------------------------------------------\n");   
     
// Write IMEM from File
write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq_ntt_inv_indirect_falcon-1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- IMEM\n");
// Read IMEM  
for (int i=0 ; i<129 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end     

 // Write DMEM from File
write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq_ntt_inv_indirect_falcon-1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- DMEM\n");
// Read DMEM  
for (int i=0 ; i<16 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end   
	   
$fwrite(f,"----------------------------------------------------------------\n");   

// Set Instruction Counter to zero (optional)
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );

// Start Programm in IMEM
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(CmdExecute), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
cc_start = cc;
// Poll on Status Register until Programm is finished
rdbk = '1;
while (rdbk != '0) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
end 

// Measure CC
cc_stop = cc; 
cc_count_falcon1024_inv_indirect = cc_stop - cc_start;        
       
// Read DMEM  
for (int i=0 ; i<1024 ; i++) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+192), .tl_o(tl_o), .tl_i(tl_i_d) );
    
    case(i)
	0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2   :   assert (rdbk == 32'd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3   :   assert (rdbk == 32'd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	5   :   assert (rdbk == 32'd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	6   :   assert (rdbk == 32'd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	7   :   assert (rdbk == 32'd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	8   :   assert (rdbk == 32'd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	9   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	10   :   assert (rdbk == 32'd10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	11   :   assert (rdbk == 32'd11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	12   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	13   :   assert (rdbk == 32'd13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	14   :   assert (rdbk == 32'd14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	15   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	16   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	17   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	18   :   assert (rdbk == 32'd18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	19   :   assert (rdbk == 32'd19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	20   :   assert (rdbk == 32'd20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	21   :   assert (rdbk == 32'd21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	22   :   assert (rdbk == 32'd22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	23   :   assert (rdbk == 32'd23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	24   :   assert (rdbk == 32'd24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	25   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	26   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	27   :   assert (rdbk == 32'd27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	28   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	29   :   assert (rdbk == 32'd29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	30   :   assert (rdbk == 32'd30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	31   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	32   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	33   :   assert (rdbk == 32'd33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	34   :   assert (rdbk == 32'd34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	35   :   assert (rdbk == 32'd35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	36   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	37   :   assert (rdbk == 32'd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	38   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	39   :   assert (rdbk == 32'd39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	40   :   assert (rdbk == 32'd40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	41   :   assert (rdbk == 32'd41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	42   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	43   :   assert (rdbk == 32'd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	44   :   assert (rdbk == 32'd44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	45   :   assert (rdbk == 32'd45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	46   :   assert (rdbk == 32'd46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	47   :   assert (rdbk == 32'd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	48   :   assert (rdbk == 32'd48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	49   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	50   :   assert (rdbk == 32'd50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	51   :   assert (rdbk == 32'd51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	52   :   assert (rdbk == 32'd52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	53   :   assert (rdbk == 32'd53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	54   :   assert (rdbk == 32'd54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	55   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	56   :   assert (rdbk == 32'd56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	57   :   assert (rdbk == 32'd57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	58   :   assert (rdbk == 32'd58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	59   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	60   :   assert (rdbk == 32'd60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	61   :   assert (rdbk == 32'd61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	62   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	63   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	64   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	65   :   assert (rdbk == 32'd65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	66   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	67   :   assert (rdbk == 32'd67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	68   :   assert (rdbk == 32'd68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	69   :   assert (rdbk == 32'd69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	70   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	71   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	72   :   assert (rdbk == 32'd72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	73   :   assert (rdbk == 32'd73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	74   :   assert (rdbk == 32'd74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	75   :   assert (rdbk == 32'd75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	76   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	77   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	78   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	79   :   assert (rdbk == 32'd79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	80   :   assert (rdbk == 32'd80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	81   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	82   :   assert (rdbk == 32'd82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	83   :   assert (rdbk == 32'd83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	84   :   assert (rdbk == 32'd84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	85   :   assert (rdbk == 32'd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	86   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	87   :   assert (rdbk == 32'd87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	88   :   assert (rdbk == 32'd88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	89   :   assert (rdbk == 32'd89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	90   :   assert (rdbk == 32'd90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	91   :   assert (rdbk == 32'd91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	92   :   assert (rdbk == 32'd92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	93   :   assert (rdbk == 32'd93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	94   :   assert (rdbk == 32'd94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	95   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	96   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	97   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	98   :   assert (rdbk == 32'd98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	99   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	100   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	101   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	102   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	103   :   assert (rdbk == 32'd103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	104   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	105   :   assert (rdbk == 32'd105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	106   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	107   :   assert (rdbk == 32'd107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	108   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	109   :   assert (rdbk == 32'd109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	110   :   assert (rdbk == 32'd110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	111   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	112   :   assert (rdbk == 32'd112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	113   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	114   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	115   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	116   :   assert (rdbk == 32'd116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	117   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	118   :   assert (rdbk == 32'd118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	119   :   assert (rdbk == 32'd119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	120   :   assert (rdbk == 32'd120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	121   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	122   :   assert (rdbk == 32'd122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	123   :   assert (rdbk == 32'd123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	124   :   assert (rdbk == 32'd124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	125   :   assert (rdbk == 32'd125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	126   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	127   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	128   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	129   :   assert (rdbk == 32'd129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	130   :   assert (rdbk == 32'd130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	131   :   assert (rdbk == 32'd131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	132   :   assert (rdbk == 32'd132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	133   :   assert (rdbk == 32'd133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	134   :   assert (rdbk == 32'd134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	135   :   assert (rdbk == 32'd135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	136   :   assert (rdbk == 32'd136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	137   :   assert (rdbk == 32'd137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	138   :   assert (rdbk == 32'd138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	139   :   assert (rdbk == 32'd139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	140   :   assert (rdbk == 32'd140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	141   :   assert (rdbk == 32'd141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	142   :   assert (rdbk == 32'd142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	143   :   assert (rdbk == 32'd143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	144   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	145   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	146   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	147   :   assert (rdbk == 32'd147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	148   :   assert (rdbk == 32'd148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	149   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	150   :   assert (rdbk == 32'd150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	151   :   assert (rdbk == 32'd151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	152   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	153   :   assert (rdbk == 32'd153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	154   :   assert (rdbk == 32'd154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	155   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	156   :   assert (rdbk == 32'd156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	157   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	158   :   assert (rdbk == 32'd158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	159   :   assert (rdbk == 32'd159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	160   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	161   :   assert (rdbk == 32'd161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	162   :   assert (rdbk == 32'd162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	163   :   assert (rdbk == 32'd163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	164   :   assert (rdbk == 32'd164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	165   :   assert (rdbk == 32'd165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	166   :   assert (rdbk == 32'd166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	167   :   assert (rdbk == 32'd167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	168   :   assert (rdbk == 32'd168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	169   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	170   :   assert (rdbk == 32'd170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	171   :   assert (rdbk == 32'd171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	172   :   assert (rdbk == 32'd172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	173   :   assert (rdbk == 32'd173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	174   :   assert (rdbk == 32'd174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	175   :   assert (rdbk == 32'd175) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	176   :   assert (rdbk == 32'd176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	177   :   assert (rdbk == 32'd177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	178   :   assert (rdbk == 32'd178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	179   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	180   :   assert (rdbk == 32'd180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	181   :   assert (rdbk == 32'd181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	182   :   assert (rdbk == 32'd182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	183   :   assert (rdbk == 32'd183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	184   :   assert (rdbk == 32'd184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	185   :   assert (rdbk == 32'd185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	186   :   assert (rdbk == 32'd186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	187   :   assert (rdbk == 32'd187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	188   :   assert (rdbk == 32'd188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	189   :   assert (rdbk == 32'd189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	190   :   assert (rdbk == 32'd190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	191   :   assert (rdbk == 32'd191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	192   :   assert (rdbk == 32'd192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	193   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	194   :   assert (rdbk == 32'd194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	195   :   assert (rdbk == 32'd195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	196   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	197   :   assert (rdbk == 32'd197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	198   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	199   :   assert (rdbk == 32'd199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	200   :   assert (rdbk == 32'd200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	201   :   assert (rdbk == 32'd201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	202   :   assert (rdbk == 32'd202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	203   :   assert (rdbk == 32'd203) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	204   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	205   :   assert (rdbk == 32'd205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	206   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	207   :   assert (rdbk == 32'd207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	208   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	209   :   assert (rdbk == 32'd209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	210   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	211   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	212   :   assert (rdbk == 32'd212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	213   :   assert (rdbk == 32'd213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	214   :   assert (rdbk == 32'd214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	215   :   assert (rdbk == 32'd215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	216   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	217   :   assert (rdbk == 32'd217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	218   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	219   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	220   :   assert (rdbk == 32'd220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	221   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	222   :   assert (rdbk == 32'd222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	223   :   assert (rdbk == 32'd223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	224   :   assert (rdbk == 32'd224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	225   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	226   :   assert (rdbk == 32'd226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	227   :   assert (rdbk == 32'd227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	228   :   assert (rdbk == 32'd228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	229   :   assert (rdbk == 32'd229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	230   :   assert (rdbk == 32'd230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	231   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	232   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	233   :   assert (rdbk == 32'd233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	234   :   assert (rdbk == 32'd234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	235   :   assert (rdbk == 32'd235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	236   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	237   :   assert (rdbk == 32'd237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	238   :   assert (rdbk == 32'd238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	239   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	240   :   assert (rdbk == 32'd240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	241   :   assert (rdbk == 32'd241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	242   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	243   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	244   :   assert (rdbk == 32'd244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	245   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	246   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	247   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	248   :   assert (rdbk == 32'd248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	249   :   assert (rdbk == 32'd249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	250   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	251   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	252   :   assert (rdbk == 32'd252) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	253   :   assert (rdbk == 32'd253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	254   :   assert (rdbk == 32'd254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	255   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	256   :   assert (rdbk == 32'd256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	257   :   assert (rdbk == 32'd257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	258   :   assert (rdbk == 32'd258) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	259   :   assert (rdbk == 32'd259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	260   :   assert (rdbk == 32'd260) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	261   :   assert (rdbk == 32'd261) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	262   :   assert (rdbk == 32'd262) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	263   :   assert (rdbk == 32'd263) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	264   :   assert (rdbk == 32'd264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	265   :   assert (rdbk == 32'd265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	266   :   assert (rdbk == 32'd266) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	267   :   assert (rdbk == 32'd267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	268   :   assert (rdbk == 32'd268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	269   :   assert (rdbk == 32'd269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	270   :   assert (rdbk == 32'd270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	271   :   assert (rdbk == 32'd271) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	272   :   assert (rdbk == 32'd272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	273   :   assert (rdbk == 32'd273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	274   :   assert (rdbk == 32'd274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	275   :   assert (rdbk == 32'd275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	276   :   assert (rdbk == 32'd276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	277   :   assert (rdbk == 32'd277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	278   :   assert (rdbk == 32'd278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	279   :   assert (rdbk == 32'd279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	280   :   assert (rdbk == 32'd280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	281   :   assert (rdbk == 32'd281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	282   :   assert (rdbk == 32'd282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	283   :   assert (rdbk == 32'd283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	284   :   assert (rdbk == 32'd284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	285   :   assert (rdbk == 32'd285) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	286   :   assert (rdbk == 32'd286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	287   :   assert (rdbk == 32'd287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	288   :   assert (rdbk == 32'd288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	289   :   assert (rdbk == 32'd289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	290   :   assert (rdbk == 32'd290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	291   :   assert (rdbk == 32'd291) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	292   :   assert (rdbk == 32'd292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	293   :   assert (rdbk == 32'd293) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	294   :   assert (rdbk == 32'd294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	295   :   assert (rdbk == 32'd295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	296   :   assert (rdbk == 32'd296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	297   :   assert (rdbk == 32'd297) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	298   :   assert (rdbk == 32'd298) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	299   :   assert (rdbk == 32'd299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	300   :   assert (rdbk == 32'd300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	301   :   assert (rdbk == 32'd301) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	302   :   assert (rdbk == 32'd302) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	303   :   assert (rdbk == 32'd303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	304   :   assert (rdbk == 32'd304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	305   :   assert (rdbk == 32'd305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	306   :   assert (rdbk == 32'd306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	307   :   assert (rdbk == 32'd307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	308   :   assert (rdbk == 32'd308) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	309   :   assert (rdbk == 32'd309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	310   :   assert (rdbk == 32'd310) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	311   :   assert (rdbk == 32'd311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	312   :   assert (rdbk == 32'd312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	313   :   assert (rdbk == 32'd313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	314   :   assert (rdbk == 32'd314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	315   :   assert (rdbk == 32'd315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	316   :   assert (rdbk == 32'd316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	317   :   assert (rdbk == 32'd317) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	318   :   assert (rdbk == 32'd318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	319   :   assert (rdbk == 32'd319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	320   :   assert (rdbk == 32'd320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	321   :   assert (rdbk == 32'd321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	322   :   assert (rdbk == 32'd322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	323   :   assert (rdbk == 32'd323) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	324   :   assert (rdbk == 32'd324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	325   :   assert (rdbk == 32'd325) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	326   :   assert (rdbk == 32'd326) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	327   :   assert (rdbk == 32'd327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	328   :   assert (rdbk == 32'd328) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	329   :   assert (rdbk == 32'd329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	330   :   assert (rdbk == 32'd330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	331   :   assert (rdbk == 32'd331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	332   :   assert (rdbk == 32'd332) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	333   :   assert (rdbk == 32'd333) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	334   :   assert (rdbk == 32'd334) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	335   :   assert (rdbk == 32'd335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	336   :   assert (rdbk == 32'd336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	337   :   assert (rdbk == 32'd337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	338   :   assert (rdbk == 32'd338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	339   :   assert (rdbk == 32'd339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	340   :   assert (rdbk == 32'd340) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	341   :   assert (rdbk == 32'd341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	342   :   assert (rdbk == 32'd342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	343   :   assert (rdbk == 32'd343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	344   :   assert (rdbk == 32'd344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	345   :   assert (rdbk == 32'd345) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	346   :   assert (rdbk == 32'd346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	347   :   assert (rdbk == 32'd347) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	348   :   assert (rdbk == 32'd348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	349   :   assert (rdbk == 32'd349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	350   :   assert (rdbk == 32'd350) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	351   :   assert (rdbk == 32'd351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	352   :   assert (rdbk == 32'd352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	353   :   assert (rdbk == 32'd353) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	354   :   assert (rdbk == 32'd354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	355   :   assert (rdbk == 32'd355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	356   :   assert (rdbk == 32'd356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	357   :   assert (rdbk == 32'd357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	358   :   assert (rdbk == 32'd358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	359   :   assert (rdbk == 32'd359) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	360   :   assert (rdbk == 32'd360) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	361   :   assert (rdbk == 32'd361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	362   :   assert (rdbk == 32'd362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	363   :   assert (rdbk == 32'd363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	364   :   assert (rdbk == 32'd364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	365   :   assert (rdbk == 32'd365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	366   :   assert (rdbk == 32'd366) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	367   :   assert (rdbk == 32'd367) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	368   :   assert (rdbk == 32'd368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	369   :   assert (rdbk == 32'd369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	370   :   assert (rdbk == 32'd370) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	371   :   assert (rdbk == 32'd371) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	372   :   assert (rdbk == 32'd372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	373   :   assert (rdbk == 32'd373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	374   :   assert (rdbk == 32'd374) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	375   :   assert (rdbk == 32'd375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	376   :   assert (rdbk == 32'd376) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	377   :   assert (rdbk == 32'd377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	378   :   assert (rdbk == 32'd378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	379   :   assert (rdbk == 32'd379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	380   :   assert (rdbk == 32'd380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	381   :   assert (rdbk == 32'd381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	382   :   assert (rdbk == 32'd382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	383   :   assert (rdbk == 32'd383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	384   :   assert (rdbk == 32'd384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	385   :   assert (rdbk == 32'd385) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	386   :   assert (rdbk == 32'd386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	387   :   assert (rdbk == 32'd387) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	388   :   assert (rdbk == 32'd388) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	389   :   assert (rdbk == 32'd389) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	390   :   assert (rdbk == 32'd390) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	391   :   assert (rdbk == 32'd391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	392   :   assert (rdbk == 32'd392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	393   :   assert (rdbk == 32'd393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	394   :   assert (rdbk == 32'd394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	395   :   assert (rdbk == 32'd395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	396   :   assert (rdbk == 32'd396) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	397   :   assert (rdbk == 32'd397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	398   :   assert (rdbk == 32'd398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	399   :   assert (rdbk == 32'd399) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	400   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	401   :   assert (rdbk == 32'd401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	402   :   assert (rdbk == 32'd402) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	403   :   assert (rdbk == 32'd403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	404   :   assert (rdbk == 32'd404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	405   :   assert (rdbk == 32'd405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	406   :   assert (rdbk == 32'd406) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	407   :   assert (rdbk == 32'd407) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	408   :   assert (rdbk == 32'd408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	409   :   assert (rdbk == 32'd409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	410   :   assert (rdbk == 32'd410) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	411   :   assert (rdbk == 32'd411) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	412   :   assert (rdbk == 32'd412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	413   :   assert (rdbk == 32'd413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	414   :   assert (rdbk == 32'd414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	415   :   assert (rdbk == 32'd415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	416   :   assert (rdbk == 32'd416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	417   :   assert (rdbk == 32'd417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	418   :   assert (rdbk == 32'd418) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	419   :   assert (rdbk == 32'd419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	420   :   assert (rdbk == 32'd420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	421   :   assert (rdbk == 32'd421) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	422   :   assert (rdbk == 32'd422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	423   :   assert (rdbk == 32'd423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	424   :   assert (rdbk == 32'd424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	425   :   assert (rdbk == 32'd425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	426   :   assert (rdbk == 32'd426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	427   :   assert (rdbk == 32'd427) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	428   :   assert (rdbk == 32'd428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	429   :   assert (rdbk == 32'd429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	430   :   assert (rdbk == 32'd430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	431   :   assert (rdbk == 32'd431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	432   :   assert (rdbk == 32'd432) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	433   :   assert (rdbk == 32'd433) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	434   :   assert (rdbk == 32'd434) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	435   :   assert (rdbk == 32'd435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	436   :   assert (rdbk == 32'd436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	437   :   assert (rdbk == 32'd437) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	438   :   assert (rdbk == 32'd438) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	439   :   assert (rdbk == 32'd439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	440   :   assert (rdbk == 32'd440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	441   :   assert (rdbk == 32'd441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	442   :   assert (rdbk == 32'd442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	443   :   assert (rdbk == 32'd443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	444   :   assert (rdbk == 32'd444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	445   :   assert (rdbk == 32'd445) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	446   :   assert (rdbk == 32'd446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	447   :   assert (rdbk == 32'd447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	448   :   assert (rdbk == 32'd448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	449   :   assert (rdbk == 32'd449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	450   :   assert (rdbk == 32'd450) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	451   :   assert (rdbk == 32'd451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	452   :   assert (rdbk == 32'd452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	453   :   assert (rdbk == 32'd453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	454   :   assert (rdbk == 32'd454) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	455   :   assert (rdbk == 32'd455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	456   :   assert (rdbk == 32'd456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	457   :   assert (rdbk == 32'd457) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	458   :   assert (rdbk == 32'd458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	459   :   assert (rdbk == 32'd459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	460   :   assert (rdbk == 32'd460) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	461   :   assert (rdbk == 32'd461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	462   :   assert (rdbk == 32'd462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	463   :   assert (rdbk == 32'd463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	464   :   assert (rdbk == 32'd464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	465   :   assert (rdbk == 32'd465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	466   :   assert (rdbk == 32'd466) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	467   :   assert (rdbk == 32'd467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	468   :   assert (rdbk == 32'd468) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	469   :   assert (rdbk == 32'd469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	470   :   assert (rdbk == 32'd470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	471   :   assert (rdbk == 32'd471) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	472   :   assert (rdbk == 32'd472) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	473   :   assert (rdbk == 32'd473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	474   :   assert (rdbk == 32'd474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	475   :   assert (rdbk == 32'd475) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	476   :   assert (rdbk == 32'd476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	477   :   assert (rdbk == 32'd477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	478   :   assert (rdbk == 32'd478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	479   :   assert (rdbk == 32'd479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	480   :   assert (rdbk == 32'd480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	481   :   assert (rdbk == 32'd481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	482   :   assert (rdbk == 32'd482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	483   :   assert (rdbk == 32'd483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	484   :   assert (rdbk == 32'd484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	485   :   assert (rdbk == 32'd485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	486   :   assert (rdbk == 32'd486) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	487   :   assert (rdbk == 32'd487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	488   :   assert (rdbk == 32'd488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	489   :   assert (rdbk == 32'd489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	490   :   assert (rdbk == 32'd490) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	491   :   assert (rdbk == 32'd491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	492   :   assert (rdbk == 32'd492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	493   :   assert (rdbk == 32'd493) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	494   :   assert (rdbk == 32'd494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	495   :   assert (rdbk == 32'd495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	496   :   assert (rdbk == 32'd496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	497   :   assert (rdbk == 32'd497) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	498   :   assert (rdbk == 32'd498) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	499   :   assert (rdbk == 32'd499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	500   :   assert (rdbk == 32'd500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	501   :   assert (rdbk == 32'd501) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	502   :   assert (rdbk == 32'd502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	503   :   assert (rdbk == 32'd503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	504   :   assert (rdbk == 32'd504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	505   :   assert (rdbk == 32'd505) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	506   :   assert (rdbk == 32'd506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	507   :   assert (rdbk == 32'd507) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	508   :   assert (rdbk == 32'd508) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	509   :   assert (rdbk == 32'd509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	510   :   assert (rdbk == 32'd510) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	511   :   assert (rdbk == 32'd511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	512   :   assert (rdbk == 32'd512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	513   :   assert (rdbk == 32'd513) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	514   :   assert (rdbk == 32'd514) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	515   :   assert (rdbk == 32'd515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	516   :   assert (rdbk == 32'd516) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	517   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	518   :   assert (rdbk == 32'd518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	519   :   assert (rdbk == 32'd519) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	520   :   assert (rdbk == 32'd520) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	521   :   assert (rdbk == 32'd521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	522   :   assert (rdbk == 32'd522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	523   :   assert (rdbk == 32'd523) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	524   :   assert (rdbk == 32'd524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	525   :   assert (rdbk == 32'd525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	526   :   assert (rdbk == 32'd526) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	527   :   assert (rdbk == 32'd527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	528   :   assert (rdbk == 32'd528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	529   :   assert (rdbk == 32'd529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	530   :   assert (rdbk == 32'd530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	531   :   assert (rdbk == 32'd531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	532   :   assert (rdbk == 32'd532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	533   :   assert (rdbk == 32'd533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	534   :   assert (rdbk == 32'd534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	535   :   assert (rdbk == 32'd535) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	536   :   assert (rdbk == 32'd536) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	537   :   assert (rdbk == 32'd537) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	538   :   assert (rdbk == 32'd538) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	539   :   assert (rdbk == 32'd539) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	540   :   assert (rdbk == 32'd540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	541   :   assert (rdbk == 32'd541) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	542   :   assert (rdbk == 32'd542) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	543   :   assert (rdbk == 32'd543) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	544   :   assert (rdbk == 32'd544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	545   :   assert (rdbk == 32'd545) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	546   :   assert (rdbk == 32'd546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	547   :   assert (rdbk == 32'd547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	548   :   assert (rdbk == 32'd548) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	549   :   assert (rdbk == 32'd549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	550   :   assert (rdbk == 32'd550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	551   :   assert (rdbk == 32'd551) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	552   :   assert (rdbk == 32'd552) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	553   :   assert (rdbk == 32'd553) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	554   :   assert (rdbk == 32'd554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	555   :   assert (rdbk == 32'd555) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	556   :   assert (rdbk == 32'd556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	557   :   assert (rdbk == 32'd557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	558   :   assert (rdbk == 32'd558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	559   :   assert (rdbk == 32'd559) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	560   :   assert (rdbk == 32'd560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	561   :   assert (rdbk == 32'd561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	562   :   assert (rdbk == 32'd562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	563   :   assert (rdbk == 32'd563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	564   :   assert (rdbk == 32'd564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	565   :   assert (rdbk == 32'd565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	566   :   assert (rdbk == 32'd566) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	567   :   assert (rdbk == 32'd567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	568   :   assert (rdbk == 32'd568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	569   :   assert (rdbk == 32'd569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	570   :   assert (rdbk == 32'd570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	571   :   assert (rdbk == 32'd571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	572   :   assert (rdbk == 32'd572) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	573   :   assert (rdbk == 32'd573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	574   :   assert (rdbk == 32'd574) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	575   :   assert (rdbk == 32'd575) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	576   :   assert (rdbk == 32'd576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	577   :   assert (rdbk == 32'd577) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	578   :   assert (rdbk == 32'd578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	579   :   assert (rdbk == 32'd579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	580   :   assert (rdbk == 32'd580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	581   :   assert (rdbk == 32'd581) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	582   :   assert (rdbk == 32'd582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	583   :   assert (rdbk == 32'd583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	584   :   assert (rdbk == 32'd584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	585   :   assert (rdbk == 32'd585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	586   :   assert (rdbk == 32'd586) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	587   :   assert (rdbk == 32'd587) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	588   :   assert (rdbk == 32'd588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	589   :   assert (rdbk == 32'd589) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	590   :   assert (rdbk == 32'd590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	591   :   assert (rdbk == 32'd591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	592   :   assert (rdbk == 32'd592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	593   :   assert (rdbk == 32'd593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	594   :   assert (rdbk == 32'd594) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	595   :   assert (rdbk == 32'd595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	596   :   assert (rdbk == 32'd596) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	597   :   assert (rdbk == 32'd597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	598   :   assert (rdbk == 32'd598) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	599   :   assert (rdbk == 32'd599) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	600   :   assert (rdbk == 32'd600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	601   :   assert (rdbk == 32'd601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	602   :   assert (rdbk == 32'd602) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	603   :   assert (rdbk == 32'd603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	604   :   assert (rdbk == 32'd604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	605   :   assert (rdbk == 32'd605) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	606   :   assert (rdbk == 32'd606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	607   :   assert (rdbk == 32'd607) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	608   :   assert (rdbk == 32'd608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	609   :   assert (rdbk == 32'd609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	610   :   assert (rdbk == 32'd610) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	611   :   assert (rdbk == 32'd611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	612   :   assert (rdbk == 32'd612) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	613   :   assert (rdbk == 32'd613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	614   :   assert (rdbk == 32'd614) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	615   :   assert (rdbk == 32'd615) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	616   :   assert (rdbk == 32'd616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	617   :   assert (rdbk == 32'd617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	618   :   assert (rdbk == 32'd618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	619   :   assert (rdbk == 32'd619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	620   :   assert (rdbk == 32'd620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	621   :   assert (rdbk == 32'd621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	622   :   assert (rdbk == 32'd622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	623   :   assert (rdbk == 32'd623) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	624   :   assert (rdbk == 32'd624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	625   :   assert (rdbk == 32'd625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	626   :   assert (rdbk == 32'd626) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	627   :   assert (rdbk == 32'd627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	628   :   assert (rdbk == 32'd628) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	629   :   assert (rdbk == 32'd629) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	630   :   assert (rdbk == 32'd630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	631   :   assert (rdbk == 32'd631) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	632   :   assert (rdbk == 32'd632) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	633   :   assert (rdbk == 32'd633) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	634   :   assert (rdbk == 32'd634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	635   :   assert (rdbk == 32'd635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	636   :   assert (rdbk == 32'd636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	637   :   assert (rdbk == 32'd637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	638   :   assert (rdbk == 32'd638) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	639   :   assert (rdbk == 32'd639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	640   :   assert (rdbk == 32'd640) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	641   :   assert (rdbk == 32'd641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	642   :   assert (rdbk == 32'd642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	643   :   assert (rdbk == 32'd643) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	644   :   assert (rdbk == 32'd644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	645   :   assert (rdbk == 32'd645) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	646   :   assert (rdbk == 32'd646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	647   :   assert (rdbk == 32'd647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	648   :   assert (rdbk == 32'd648) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	649   :   assert (rdbk == 32'd649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	650   :   assert (rdbk == 32'd650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	651   :   assert (rdbk == 32'd651) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	652   :   assert (rdbk == 32'd652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	653   :   assert (rdbk == 32'd653) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	654   :   assert (rdbk == 32'd654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	655   :   assert (rdbk == 32'd655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	656   :   assert (rdbk == 32'd656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	657   :   assert (rdbk == 32'd657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	658   :   assert (rdbk == 32'd658) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	659   :   assert (rdbk == 32'd659) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	660   :   assert (rdbk == 32'd660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	661   :   assert (rdbk == 32'd661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	662   :   assert (rdbk == 32'd662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	663   :   assert (rdbk == 32'd663) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	664   :   assert (rdbk == 32'd664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	665   :   assert (rdbk == 32'd665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	666   :   assert (rdbk == 32'd666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	667   :   assert (rdbk == 32'd667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	668   :   assert (rdbk == 32'd668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	669   :   assert (rdbk == 32'd669) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	670   :   assert (rdbk == 32'd670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	671   :   assert (rdbk == 32'd671) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	672   :   assert (rdbk == 32'd672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	673   :   assert (rdbk == 32'd673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	674   :   assert (rdbk == 32'd674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	675   :   assert (rdbk == 32'd675) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	676   :   assert (rdbk == 32'd676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	677   :   assert (rdbk == 32'd677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	678   :   assert (rdbk == 32'd678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	679   :   assert (rdbk == 32'd679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	680   :   assert (rdbk == 32'd680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	681   :   assert (rdbk == 32'd681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	682   :   assert (rdbk == 32'd682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	683   :   assert (rdbk == 32'd683) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	684   :   assert (rdbk == 32'd684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	685   :   assert (rdbk == 32'd685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	686   :   assert (rdbk == 32'd686) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	687   :   assert (rdbk == 32'd687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	688   :   assert (rdbk == 32'd688) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	689   :   assert (rdbk == 32'd689) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	690   :   assert (rdbk == 32'd690) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	691   :   assert (rdbk == 32'd691) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	692   :   assert (rdbk == 32'd692) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	693   :   assert (rdbk == 32'd693) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	694   :   assert (rdbk == 32'd694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	695   :   assert (rdbk == 32'd695) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	696   :   assert (rdbk == 32'd696) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	697   :   assert (rdbk == 32'd697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	698   :   assert (rdbk == 32'd698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	699   :   assert (rdbk == 32'd699) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	700   :   assert (rdbk == 32'd700) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	701   :   assert (rdbk == 32'd701) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	702   :   assert (rdbk == 32'd702) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	703   :   assert (rdbk == 32'd703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	704   :   assert (rdbk == 32'd704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	705   :   assert (rdbk == 32'd705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	706   :   assert (rdbk == 32'd706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	707   :   assert (rdbk == 32'd707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	708   :   assert (rdbk == 32'd708) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	709   :   assert (rdbk == 32'd709) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	710   :   assert (rdbk == 32'd710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	711   :   assert (rdbk == 32'd711) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	712   :   assert (rdbk == 32'd712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	713   :   assert (rdbk == 32'd713) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	714   :   assert (rdbk == 32'd714) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	715   :   assert (rdbk == 32'd715) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	716   :   assert (rdbk == 32'd716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	717   :   assert (rdbk == 32'd717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	718   :   assert (rdbk == 32'd718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	719   :   assert (rdbk == 32'd719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	720   :   assert (rdbk == 32'd720) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	721   :   assert (rdbk == 32'd721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	722   :   assert (rdbk == 32'd722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	723   :   assert (rdbk == 32'd723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	724   :   assert (rdbk == 32'd724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	725   :   assert (rdbk == 32'd725) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	726   :   assert (rdbk == 32'd726) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	727   :   assert (rdbk == 32'd727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	728   :   assert (rdbk == 32'd728) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	729   :   assert (rdbk == 32'd729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	730   :   assert (rdbk == 32'd730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	731   :   assert (rdbk == 32'd731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	732   :   assert (rdbk == 32'd732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	733   :   assert (rdbk == 32'd733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	734   :   assert (rdbk == 32'd734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	735   :   assert (rdbk == 32'd735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	736   :   assert (rdbk == 32'd736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	737   :   assert (rdbk == 32'd737) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	738   :   assert (rdbk == 32'd738) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	739   :   assert (rdbk == 32'd739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	740   :   assert (rdbk == 32'd740) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	741   :   assert (rdbk == 32'd741) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	742   :   assert (rdbk == 32'd742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	743   :   assert (rdbk == 32'd743) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	744   :   assert (rdbk == 32'd744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	745   :   assert (rdbk == 32'd745) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	746   :   assert (rdbk == 32'd746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	747   :   assert (rdbk == 32'd747) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	748   :   assert (rdbk == 32'd748) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	749   :   assert (rdbk == 32'd749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	750   :   assert (rdbk == 32'd750) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	751   :   assert (rdbk == 32'd751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	752   :   assert (rdbk == 32'd752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	753   :   assert (rdbk == 32'd753) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	754   :   assert (rdbk == 32'd754) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	755   :   assert (rdbk == 32'd755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	756   :   assert (rdbk == 32'd756) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	757   :   assert (rdbk == 32'd757) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	758   :   assert (rdbk == 32'd758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	759   :   assert (rdbk == 32'd759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	760   :   assert (rdbk == 32'd760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	761   :   assert (rdbk == 32'd761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	762   :   assert (rdbk == 32'd762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	763   :   assert (rdbk == 32'd763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	764   :   assert (rdbk == 32'd764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	765   :   assert (rdbk == 32'd765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	766   :   assert (rdbk == 32'd766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	767   :   assert (rdbk == 32'd767) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	768   :   assert (rdbk == 32'd768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	769   :   assert (rdbk == 32'd769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	770   :   assert (rdbk == 32'd770) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	771   :   assert (rdbk == 32'd771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	772   :   assert (rdbk == 32'd772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	773   :   assert (rdbk == 32'd773) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	774   :   assert (rdbk == 32'd774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	775   :   assert (rdbk == 32'd775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	776   :   assert (rdbk == 32'd776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	777   :   assert (rdbk == 32'd777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	778   :   assert (rdbk == 32'd778) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	779   :   assert (rdbk == 32'd779) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	780   :   assert (rdbk == 32'd780) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	781   :   assert (rdbk == 32'd781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	782   :   assert (rdbk == 32'd782) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	783   :   assert (rdbk == 32'd783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	784   :   assert (rdbk == 32'd784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	785   :   assert (rdbk == 32'd785) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	786   :   assert (rdbk == 32'd786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	787   :   assert (rdbk == 32'd787) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	788   :   assert (rdbk == 32'd788) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	789   :   assert (rdbk == 32'd789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	790   :   assert (rdbk == 32'd790) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	791   :   assert (rdbk == 32'd791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	792   :   assert (rdbk == 32'd792) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	793   :   assert (rdbk == 32'd793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	794   :   assert (rdbk == 32'd794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	795   :   assert (rdbk == 32'd795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	796   :   assert (rdbk == 32'd796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	797   :   assert (rdbk == 32'd797) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	798   :   assert (rdbk == 32'd798) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	799   :   assert (rdbk == 32'd799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	800   :   assert (rdbk == 32'd800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	801   :   assert (rdbk == 32'd801) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	802   :   assert (rdbk == 32'd802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	803   :   assert (rdbk == 32'd803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	804   :   assert (rdbk == 32'd804) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	805   :   assert (rdbk == 32'd805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	806   :   assert (rdbk == 32'd806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	807   :   assert (rdbk == 32'd807) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	808   :   assert (rdbk == 32'd808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	809   :   assert (rdbk == 32'd809) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	810   :   assert (rdbk == 32'd810) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	811   :   assert (rdbk == 32'd811) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	812   :   assert (rdbk == 32'd812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	813   :   assert (rdbk == 32'd813) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	814   :   assert (rdbk == 32'd814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	815   :   assert (rdbk == 32'd815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	816   :   assert (rdbk == 32'd816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	817   :   assert (rdbk == 32'd817) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	818   :   assert (rdbk == 32'd818) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	819   :   assert (rdbk == 32'd819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	820   :   assert (rdbk == 32'd820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	821   :   assert (rdbk == 32'd821) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	822   :   assert (rdbk == 32'd822) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	823   :   assert (rdbk == 32'd823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	824   :   assert (rdbk == 32'd824) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	825   :   assert (rdbk == 32'd825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	826   :   assert (rdbk == 32'd826) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	827   :   assert (rdbk == 32'd827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	828   :   assert (rdbk == 32'd828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	829   :   assert (rdbk == 32'd829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	830   :   assert (rdbk == 32'd830) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	831   :   assert (rdbk == 32'd831) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	832   :   assert (rdbk == 32'd832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	833   :   assert (rdbk == 32'd833) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	834   :   assert (rdbk == 32'd834) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	835   :   assert (rdbk == 32'd835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	836   :   assert (rdbk == 32'd836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	837   :   assert (rdbk == 32'd837) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	838   :   assert (rdbk == 32'd838) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	839   :   assert (rdbk == 32'd839) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	840   :   assert (rdbk == 32'd840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	841   :   assert (rdbk == 32'd841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	842   :   assert (rdbk == 32'd842) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	843   :   assert (rdbk == 32'd843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	844   :   assert (rdbk == 32'd844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	845   :   assert (rdbk == 32'd845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	846   :   assert (rdbk == 32'd846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	847   :   assert (rdbk == 32'd847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	848   :   assert (rdbk == 32'd848) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	849   :   assert (rdbk == 32'd849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	850   :   assert (rdbk == 32'd850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	851   :   assert (rdbk == 32'd851) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	852   :   assert (rdbk == 32'd852) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	853   :   assert (rdbk == 32'd853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	854   :   assert (rdbk == 32'd854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	855   :   assert (rdbk == 32'd855) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	856   :   assert (rdbk == 32'd856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	857   :   assert (rdbk == 32'd857) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	858   :   assert (rdbk == 32'd858) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	859   :   assert (rdbk == 32'd859) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	860   :   assert (rdbk == 32'd860) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	861   :   assert (rdbk == 32'd861) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	862   :   assert (rdbk == 32'd862) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	863   :   assert (rdbk == 32'd863) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	864   :   assert (rdbk == 32'd864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	865   :   assert (rdbk == 32'd865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	866   :   assert (rdbk == 32'd866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	867   :   assert (rdbk == 32'd867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	868   :   assert (rdbk == 32'd868) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	869   :   assert (rdbk == 32'd869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	870   :   assert (rdbk == 32'd870) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	871   :   assert (rdbk == 32'd871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	872   :   assert (rdbk == 32'd872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	873   :   assert (rdbk == 32'd873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	874   :   assert (rdbk == 32'd874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	875   :   assert (rdbk == 32'd875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	876   :   assert (rdbk == 32'd876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	877   :   assert (rdbk == 32'd877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	878   :   assert (rdbk == 32'd878) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	879   :   assert (rdbk == 32'd879) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	880   :   assert (rdbk == 32'd880) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	881   :   assert (rdbk == 32'd881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	882   :   assert (rdbk == 32'd882) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	883   :   assert (rdbk == 32'd883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	884   :   assert (rdbk == 32'd884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	885   :   assert (rdbk == 32'd885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	886   :   assert (rdbk == 32'd886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	887   :   assert (rdbk == 32'd887) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	888   :   assert (rdbk == 32'd888) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	889   :   assert (rdbk == 32'd889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	890   :   assert (rdbk == 32'd890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	891   :   assert (rdbk == 32'd891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	892   :   assert (rdbk == 32'd892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	893   :   assert (rdbk == 32'd893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	894   :   assert (rdbk == 32'd894) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	895   :   assert (rdbk == 32'd895) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	896   :   assert (rdbk == 32'd896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	897   :   assert (rdbk == 32'd897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	898   :   assert (rdbk == 32'd898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	899   :   assert (rdbk == 32'd899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	900   :   assert (rdbk == 32'd900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	901   :   assert (rdbk == 32'd901) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	902   :   assert (rdbk == 32'd902) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	903   :   assert (rdbk == 32'd903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	904   :   assert (rdbk == 32'd904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	905   :   assert (rdbk == 32'd905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	906   :   assert (rdbk == 32'd906) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	907   :   assert (rdbk == 32'd907) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	908   :   assert (rdbk == 32'd908) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	909   :   assert (rdbk == 32'd909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	910   :   assert (rdbk == 32'd910) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	911   :   assert (rdbk == 32'd911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	912   :   assert (rdbk == 32'd912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	913   :   assert (rdbk == 32'd913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	914   :   assert (rdbk == 32'd914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	915   :   assert (rdbk == 32'd915) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	916   :   assert (rdbk == 32'd916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	917   :   assert (rdbk == 32'd917) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	918   :   assert (rdbk == 32'd918) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	919   :   assert (rdbk == 32'd919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	920   :   assert (rdbk == 32'd920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	921   :   assert (rdbk == 32'd921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	922   :   assert (rdbk == 32'd922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	923   :   assert (rdbk == 32'd923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	924   :   assert (rdbk == 32'd924) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	925   :   assert (rdbk == 32'd925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	926   :   assert (rdbk == 32'd926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	927   :   assert (rdbk == 32'd927) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	928   :   assert (rdbk == 32'd928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	929   :   assert (rdbk == 32'd929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	930   :   assert (rdbk == 32'd930) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	931   :   assert (rdbk == 32'd931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	932   :   assert (rdbk == 32'd932) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	933   :   assert (rdbk == 32'd933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	934   :   assert (rdbk == 32'd934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	935   :   assert (rdbk == 32'd935) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	936   :   assert (rdbk == 32'd936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	937   :   assert (rdbk == 32'd937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	938   :   assert (rdbk == 32'd938) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	939   :   assert (rdbk == 32'd939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	940   :   assert (rdbk == 32'd940) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	941   :   assert (rdbk == 32'd941) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	942   :   assert (rdbk == 32'd942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	943   :   assert (rdbk == 32'd943) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	944   :   assert (rdbk == 32'd944) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	945   :   assert (rdbk == 32'd945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	946   :   assert (rdbk == 32'd946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	947   :   assert (rdbk == 32'd947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	948   :   assert (rdbk == 32'd948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	949   :   assert (rdbk == 32'd949) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	950   :   assert (rdbk == 32'd950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	951   :   assert (rdbk == 32'd951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	952   :   assert (rdbk == 32'd952) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	953   :   assert (rdbk == 32'd953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	954   :   assert (rdbk == 32'd954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	955   :   assert (rdbk == 32'd955) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	956   :   assert (rdbk == 32'd956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	957   :   assert (rdbk == 32'd957) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	958   :   assert (rdbk == 32'd958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	959   :   assert (rdbk == 32'd959) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	960   :   assert (rdbk == 32'd960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	961   :   assert (rdbk == 32'd961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	962   :   assert (rdbk == 32'd962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	963   :   assert (rdbk == 32'd963) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	964   :   assert (rdbk == 32'd964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	965   :   assert (rdbk == 32'd965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	966   :   assert (rdbk == 32'd966) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	967   :   assert (rdbk == 32'd967) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	968   :   assert (rdbk == 32'd968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	969   :   assert (rdbk == 32'd969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	970   :   assert (rdbk == 32'd970) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	971   :   assert (rdbk == 32'd971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	972   :   assert (rdbk == 32'd972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	973   :   assert (rdbk == 32'd973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	974   :   assert (rdbk == 32'd974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	975   :   assert (rdbk == 32'd975) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	976   :   assert (rdbk == 32'd976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	977   :   assert (rdbk == 32'd977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	978   :   assert (rdbk == 32'd978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	979   :   assert (rdbk == 32'd979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	980   :   assert (rdbk == 32'd980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	981   :   assert (rdbk == 32'd981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	982   :   assert (rdbk == 32'd982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	983   :   assert (rdbk == 32'd983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	984   :   assert (rdbk == 32'd984) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	985   :   assert (rdbk == 32'd985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	986   :   assert (rdbk == 32'd986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	987   :   assert (rdbk == 32'd987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	988   :   assert (rdbk == 32'd988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	989   :   assert (rdbk == 32'd989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	990   :   assert (rdbk == 32'd990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	991   :   assert (rdbk == 32'd991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	992   :   assert (rdbk == 32'd992) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	993   :   assert (rdbk == 32'd993) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	994   :   assert (rdbk == 32'd994) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	995   :   assert (rdbk == 32'd995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	996   :   assert (rdbk == 32'd996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	997   :   assert (rdbk == 32'd997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	998   :   assert (rdbk == 32'd998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	999   :   assert (rdbk == 32'd999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1000   :   assert (rdbk == 32'd1000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1001   :   assert (rdbk == 32'd1001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1002   :   assert (rdbk == 32'd1002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1003   :   assert (rdbk == 32'd1003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1004   :   assert (rdbk == 32'd1004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1005   :   assert (rdbk == 32'd1005) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1006   :   assert (rdbk == 32'd1006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1007   :   assert (rdbk == 32'd1007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1008   :   assert (rdbk == 32'd1008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1009   :   assert (rdbk == 32'd1009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1010   :   assert (rdbk == 32'd1010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1011   :   assert (rdbk == 32'd1011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1012   :   assert (rdbk == 32'd1012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1013   :   assert (rdbk == 32'd1013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1014   :   assert (rdbk == 32'd1014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1015   :   assert (rdbk == 32'd1015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1016   :   assert (rdbk == 32'd1016) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1017   :   assert (rdbk == 32'd1017) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1018   :   assert (rdbk == 32'd1018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1019   :   assert (rdbk == 32'd1019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1020   :   assert (rdbk == 32'd1020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1021   :   assert (rdbk == 32'd1021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1022   :   assert (rdbk == 32'd1022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1023   :   assert (rdbk == 32'd1023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
    endcase
end

