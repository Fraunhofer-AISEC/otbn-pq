// Copyright Copyright Fraunhofer Institute for Applied and Integrated Security (AISEC).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

$fwrite(f,"----------------------------------------------------------------\n");   
$fwrite(f,"-- PQ-NTT-Indirect (Falcon-512)\n");
$fwrite(f,"----------------------------------------------------------------\n");   
     
// Write IMEM from File
write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq_ntt_indirect_falcon-512.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- IMEM\n");
// Read IMEM  
for (int i=0 ; i<129 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end     

 // Write DMEM from File
write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq_ntt_indirect_falcon-512.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- DMEM\n");
// Read DMEM  
for (int i=0 ; i<16 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end   
	   
$fwrite(f,"----------------------------------------------------------------\n");   

// Set Instruction Counter to zero (optional)
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );

// Start Programm in IMEM
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(CmdExecute), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
cc_start = cc;
// Poll on Status Register until Programm is finished
rdbk = '1;
while (rdbk != '0) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
end 

// Measure CC
cc_stop = cc; 
cc_count_falcon512_indirect = cc_stop - cc_start;        
       
// Read DMEM  
for (int i=0 ; i<512 ; i++) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+192), .tl_o(tl_o), .tl_i(tl_i_d) );
    
    case(i)
	0   :   assert (rdbk == 32'd3478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1   :   assert (rdbk == 32'd8305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2   :   assert (rdbk == 32'd9294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3   :   assert (rdbk == 32'd9394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4   :   assert (rdbk == 32'd6662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	5   :   assert (rdbk == 32'd5985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	6   :   assert (rdbk == 32'd3132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	7   :   assert (rdbk == 32'd5560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	8   :   assert (rdbk == 32'd8657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	9   :   assert (rdbk == 32'd3644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	10   :   assert (rdbk == 32'd8479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	11   :   assert (rdbk == 32'd11062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	12   :   assert (rdbk == 32'd358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	13   :   assert (rdbk == 32'd10395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	14   :   assert (rdbk == 32'd9828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	15   :   assert (rdbk == 32'd11980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	16   :   assert (rdbk == 32'd6723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	17   :   assert (rdbk == 32'd365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	18   :   assert (rdbk == 32'd6206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	19   :   assert (rdbk == 32'd8244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	20   :   assert (rdbk == 32'd9116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	21   :   assert (rdbk == 32'd8799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	22   :   assert (rdbk == 32'd1938) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	23   :   assert (rdbk == 32'd6517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	24   :   assert (rdbk == 32'd3491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	25   :   assert (rdbk == 32'd8590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	26   :   assert (rdbk == 32'd4573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	27   :   assert (rdbk == 32'd3003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	28   :   assert (rdbk == 32'd8920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	29   :   assert (rdbk == 32'd6129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	30   :   assert (rdbk == 32'd1131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	31   :   assert (rdbk == 32'd3898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	32   :   assert (rdbk == 32'd6024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	33   :   assert (rdbk == 32'd4583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	34   :   assert (rdbk == 32'd1222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	35   :   assert (rdbk == 32'd2936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	36   :   assert (rdbk == 32'd8324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	37   :   assert (rdbk == 32'd12266) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	38   :   assert (rdbk == 32'd4260) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	39   :   assert (rdbk == 32'd3294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	40   :   assert (rdbk == 32'd6324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	41   :   assert (rdbk == 32'd6173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	42   :   assert (rdbk == 32'd1261) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	43   :   assert (rdbk == 32'd11311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	44   :   assert (rdbk == 32'd1985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	45   :   assert (rdbk == 32'd5436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	46   :   assert (rdbk == 32'd10597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	47   :   assert (rdbk == 32'd4052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	48   :   assert (rdbk == 32'd6793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	49   :   assert (rdbk == 32'd8528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	50   :   assert (rdbk == 32'd10528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	51   :   assert (rdbk == 32'd9185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	52   :   assert (rdbk == 32'd7661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	53   :   assert (rdbk == 32'd7160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	54   :   assert (rdbk == 32'd11694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	55   :   assert (rdbk == 32'd10504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	56   :   assert (rdbk == 32'd8452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	57   :   assert (rdbk == 32'd5370) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	58   :   assert (rdbk == 32'd4710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	59   :   assert (rdbk == 32'd12110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	60   :   assert (rdbk == 32'd4970) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	61   :   assert (rdbk == 32'd10967) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	62   :   assert (rdbk == 32'd6398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	63   :   assert (rdbk == 32'd5014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	64   :   assert (rdbk == 32'd5208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	65   :   assert (rdbk == 32'd5550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	66   :   assert (rdbk == 32'd4549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	67   :   assert (rdbk == 32'd3126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	68   :   assert (rdbk == 32'd10965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	69   :   assert (rdbk == 32'd7128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	70   :   assert (rdbk == 32'd7412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	71   :   assert (rdbk == 32'd4171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	72   :   assert (rdbk == 32'd6892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	73   :   assert (rdbk == 32'd8806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	74   :   assert (rdbk == 32'd12189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	75   :   assert (rdbk == 32'd10672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	76   :   assert (rdbk == 32'd8860) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	77   :   assert (rdbk == 32'd11349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	78   :   assert (rdbk == 32'd10792) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	79   :   assert (rdbk == 32'd2003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	80   :   assert (rdbk == 32'd7810) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	81   :   assert (rdbk == 32'd11972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	82   :   assert (rdbk == 32'd8697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	83   :   assert (rdbk == 32'd11170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	84   :   assert (rdbk == 32'd4625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	85   :   assert (rdbk == 32'd9323) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	86   :   assert (rdbk == 32'd2483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	87   :   assert (rdbk == 32'd4636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	88   :   assert (rdbk == 32'd2111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	89   :   assert (rdbk == 32'd8997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	90   :   assert (rdbk == 32'd3674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	91   :   assert (rdbk == 32'd922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	92   :   assert (rdbk == 32'd6965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	93   :   assert (rdbk == 32'd2760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	94   :   assert (rdbk == 32'd11138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	95   :   assert (rdbk == 32'd4506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	96   :   assert (rdbk == 32'd2302) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	97   :   assert (rdbk == 32'd9304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	98   :   assert (rdbk == 32'd3880) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	99   :   assert (rdbk == 32'd5867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	100   :   assert (rdbk == 32'd3166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	101   :   assert (rdbk == 32'd6674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	102   :   assert (rdbk == 32'd6735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	103   :   assert (rdbk == 32'd5522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	104   :   assert (rdbk == 32'd5118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	105   :   assert (rdbk == 32'd8941) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	106   :   assert (rdbk == 32'd7341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	107   :   assert (rdbk == 32'd11250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	108   :   assert (rdbk == 32'd10319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	109   :   assert (rdbk == 32'd4613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	110   :   assert (rdbk == 32'd8373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	111   :   assert (rdbk == 32'd11294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	112   :   assert (rdbk == 32'd8083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	113   :   assert (rdbk == 32'd7760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	114   :   assert (rdbk == 32'd5583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	115   :   assert (rdbk == 32'd4772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	116   :   assert (rdbk == 32'd9982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	117   :   assert (rdbk == 32'd1698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	118   :   assert (rdbk == 32'd6634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	119   :   assert (rdbk == 32'd12261) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	120   :   assert (rdbk == 32'd8451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	121   :   assert (rdbk == 32'd1812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	122   :   assert (rdbk == 32'd3451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	123   :   assert (rdbk == 32'd621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	124   :   assert (rdbk == 32'd4584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	125   :   assert (rdbk == 32'd8591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	126   :   assert (rdbk == 32'd1331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	127   :   assert (rdbk == 32'd1083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	128   :   assert (rdbk == 32'd5759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	129   :   assert (rdbk == 32'd1373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	130   :   assert (rdbk == 32'd730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	131   :   assert (rdbk == 32'd7998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	132   :   assert (rdbk == 32'd2942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	133   :   assert (rdbk == 32'd10805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	134   :   assert (rdbk == 32'd5448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	135   :   assert (rdbk == 32'd953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	136   :   assert (rdbk == 32'd10679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	137   :   assert (rdbk == 32'd1256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	138   :   assert (rdbk == 32'd7046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	139   :   assert (rdbk == 32'd492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	140   :   assert (rdbk == 32'd6316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	141   :   assert (rdbk == 32'd5909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	142   :   assert (rdbk == 32'd9654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	143   :   assert (rdbk == 32'd11764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	144   :   assert (rdbk == 32'd7025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	145   :   assert (rdbk == 32'd7611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	146   :   assert (rdbk == 32'd2889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	147   :   assert (rdbk == 32'd3751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	148   :   assert (rdbk == 32'd6172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	149   :   assert (rdbk == 32'd6391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	150   :   assert (rdbk == 32'd10611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	151   :   assert (rdbk == 32'd7941) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	152   :   assert (rdbk == 32'd7563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	153   :   assert (rdbk == 32'd11079) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	154   :   assert (rdbk == 32'd4588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	155   :   assert (rdbk == 32'd10690) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	156   :   assert (rdbk == 32'd3865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	157   :   assert (rdbk == 32'd3033) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	158   :   assert (rdbk == 32'd6576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	159   :   assert (rdbk == 32'd4322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	160   :   assert (rdbk == 32'd2099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	161   :   assert (rdbk == 32'd2549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	162   :   assert (rdbk == 32'd4041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	163   :   assert (rdbk == 32'd1904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	164   :   assert (rdbk == 32'd10519) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	165   :   assert (rdbk == 32'd7012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	166   :   assert (rdbk == 32'd10196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	167   :   assert (rdbk == 32'd7732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	168   :   assert (rdbk == 32'd9827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	169   :   assert (rdbk == 32'd10792) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	170   :   assert (rdbk == 32'd4816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	171   :   assert (rdbk == 32'd9771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	172   :   assert (rdbk == 32'd590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	173   :   assert (rdbk == 32'd7304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	174   :   assert (rdbk == 32'd8031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	175   :   assert (rdbk == 32'd5521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	176   :   assert (rdbk == 32'd9032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	177   :   assert (rdbk == 32'd1620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	178   :   assert (rdbk == 32'd4101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	179   :   assert (rdbk == 32'd4303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	180   :   assert (rdbk == 32'd5499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	181   :   assert (rdbk == 32'd7620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	182   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	183   :   assert (rdbk == 32'd10736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	184   :   assert (rdbk == 32'd8642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	185   :   assert (rdbk == 32'd3430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	186   :   assert (rdbk == 32'd8118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	187   :   assert (rdbk == 32'd8166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	188   :   assert (rdbk == 32'd4877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	189   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	190   :   assert (rdbk == 32'd5304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	191   :   assert (rdbk == 32'd7964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	192   :   assert (rdbk == 32'd5063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	193   :   assert (rdbk == 32'd4584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	194   :   assert (rdbk == 32'd9487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	195   :   assert (rdbk == 32'd8348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	196   :   assert (rdbk == 32'd1734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	197   :   assert (rdbk == 32'd2939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	198   :   assert (rdbk == 32'd6958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	199   :   assert (rdbk == 32'd10013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	200   :   assert (rdbk == 32'd3391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	201   :   assert (rdbk == 32'd2562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	202   :   assert (rdbk == 32'd5609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	203   :   assert (rdbk == 32'd4459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	204   :   assert (rdbk == 32'd1997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	205   :   assert (rdbk == 32'd9743) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	206   :   assert (rdbk == 32'd5443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	207   :   assert (rdbk == 32'd10604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	208   :   assert (rdbk == 32'd8722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	209   :   assert (rdbk == 32'd8368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	210   :   assert (rdbk == 32'd6139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	211   :   assert (rdbk == 32'd1825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	212   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	213   :   assert (rdbk == 32'd5461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	214   :   assert (rdbk == 32'd2520) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	215   :   assert (rdbk == 32'd796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	216   :   assert (rdbk == 32'd8926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	217   :   assert (rdbk == 32'd11417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	218   :   assert (rdbk == 32'd9476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	219   :   assert (rdbk == 32'd5541) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	220   :   assert (rdbk == 32'd11866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	221   :   assert (rdbk == 32'd10839) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	222   :   assert (rdbk == 32'd5724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	223   :   assert (rdbk == 32'd1746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	224   :   assert (rdbk == 32'd3344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	225   :   assert (rdbk == 32'd7852) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	226   :   assert (rdbk == 32'd8762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	227   :   assert (rdbk == 32'd4351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	228   :   assert (rdbk == 32'd4068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	229   :   assert (rdbk == 32'd11749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	230   :   assert (rdbk == 32'd5791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	231   :   assert (rdbk == 32'd8103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	232   :   assert (rdbk == 32'd7939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	233   :   assert (rdbk == 32'd7956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	234   :   assert (rdbk == 32'd12126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	235   :   assert (rdbk == 32'd10206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	236   :   assert (rdbk == 32'd6319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	237   :   assert (rdbk == 32'd1253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	238   :   assert (rdbk == 32'd7230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	239   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	240   :   assert (rdbk == 32'd8230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	241   :   assert (rdbk == 32'd4957) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	242   :   assert (rdbk == 32'd5750) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	243   :   assert (rdbk == 32'd583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	244   :   assert (rdbk == 32'd3127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	245   :   assert (rdbk == 32'd5092) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	246   :   assert (rdbk == 32'd2272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	247   :   assert (rdbk == 32'd6433) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	248   :   assert (rdbk == 32'd6886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	249   :   assert (rdbk == 32'd2221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	250   :   assert (rdbk == 32'd4352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	251   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	252   :   assert (rdbk == 32'd1973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	253   :   assert (rdbk == 32'd8419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	254   :   assert (rdbk == 32'd3058) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	255   :   assert (rdbk == 32'd10731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	256   :   assert (rdbk == 32'd832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	257   :   assert (rdbk == 32'd8073) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	258   :   assert (rdbk == 32'd11453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	259   :   assert (rdbk == 32'd6766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	260   :   assert (rdbk == 32'd6306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	261   :   assert (rdbk == 32'd10507) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	262   :   assert (rdbk == 32'd9219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	263   :   assert (rdbk == 32'd4911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	264   :   assert (rdbk == 32'd320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	265   :   assert (rdbk == 32'd4352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	266   :   assert (rdbk == 32'd9126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	267   :   assert (rdbk == 32'd9699) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	268   :   assert (rdbk == 32'd3267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	269   :   assert (rdbk == 32'd10701) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	270   :   assert (rdbk == 32'd7238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	271   :   assert (rdbk == 32'd4245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	272   :   assert (rdbk == 32'd11832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	273   :   assert (rdbk == 32'd4718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	274   :   assert (rdbk == 32'd4207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	275   :   assert (rdbk == 32'd11117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	276   :   assert (rdbk == 32'd2188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	277   :   assert (rdbk == 32'd5184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	278   :   assert (rdbk == 32'd1664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	279   :   assert (rdbk == 32'd413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	280   :   assert (rdbk == 32'd3331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	281   :   assert (rdbk == 32'd9465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	282   :   assert (rdbk == 32'd6620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	283   :   assert (rdbk == 32'd3116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	284   :   assert (rdbk == 32'd5582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	285   :   assert (rdbk == 32'd3095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	286   :   assert (rdbk == 32'd9987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	287   :   assert (rdbk == 32'd9217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	288   :   assert (rdbk == 32'd673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	289   :   assert (rdbk == 32'd10393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	290   :   assert (rdbk == 32'd7383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	291   :   assert (rdbk == 32'd11335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	292   :   assert (rdbk == 32'd7057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	293   :   assert (rdbk == 32'd343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	294   :   assert (rdbk == 32'd2100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	295   :   assert (rdbk == 32'd10387) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	296   :   assert (rdbk == 32'd11657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	297   :   assert (rdbk == 32'd3197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	298   :   assert (rdbk == 32'd6384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	299   :   assert (rdbk == 32'd2256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	300   :   assert (rdbk == 32'd7195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	301   :   assert (rdbk == 32'd8966) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	302   :   assert (rdbk == 32'd6343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	303   :   assert (rdbk == 32'd9782) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	304   :   assert (rdbk == 32'd10562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	305   :   assert (rdbk == 32'd3883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	306   :   assert (rdbk == 32'd9990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	307   :   assert (rdbk == 32'd6143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	308   :   assert (rdbk == 32'd6579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	309   :   assert (rdbk == 32'd10741) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	310   :   assert (rdbk == 32'd8973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	311   :   assert (rdbk == 32'd1239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	312   :   assert (rdbk == 32'd6050) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	313   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	314   :   assert (rdbk == 32'd9572) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	315   :   assert (rdbk == 32'd6346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	316   :   assert (rdbk == 32'd10825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	317   :   assert (rdbk == 32'd6755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	318   :   assert (rdbk == 32'd3082) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	319   :   assert (rdbk == 32'd6983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	320   :   assert (rdbk == 32'd4599) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	321   :   assert (rdbk == 32'd12059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	322   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	323   :   assert (rdbk == 32'd1596) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	324   :   assert (rdbk == 32'd11382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	325   :   assert (rdbk == 32'd2269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	326   :   assert (rdbk == 32'd7426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	327   :   assert (rdbk == 32'd1130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	328   :   assert (rdbk == 32'd6312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	329   :   assert (rdbk == 32'd3563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	330   :   assert (rdbk == 32'd914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	331   :   assert (rdbk == 32'd1410) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	332   :   assert (rdbk == 32'd10019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	333   :   assert (rdbk == 32'd12179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	334   :   assert (rdbk == 32'd3443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	335   :   assert (rdbk == 32'd11670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	336   :   assert (rdbk == 32'd12005) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	337   :   assert (rdbk == 32'd1256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	338   :   assert (rdbk == 32'd1812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	339   :   assert (rdbk == 32'd4928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	340   :   assert (rdbk == 32'd299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	341   :   assert (rdbk == 32'd6449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	342   :   assert (rdbk == 32'd10435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	343   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	344   :   assert (rdbk == 32'd6703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	345   :   assert (rdbk == 32'd5618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	346   :   assert (rdbk == 32'd7229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	347   :   assert (rdbk == 32'd8046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	348   :   assert (rdbk == 32'd3908) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	349   :   assert (rdbk == 32'd3485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	350   :   assert (rdbk == 32'd9999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	351   :   assert (rdbk == 32'd8409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	352   :   assert (rdbk == 32'd5716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	353   :   assert (rdbk == 32'd9779) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	354   :   assert (rdbk == 32'd10612) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	355   :   assert (rdbk == 32'd10113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	356   :   assert (rdbk == 32'd7087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	357   :   assert (rdbk == 32'd2728) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	358   :   assert (rdbk == 32'd9673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	359   :   assert (rdbk == 32'd10156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	360   :   assert (rdbk == 32'd7131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	361   :   assert (rdbk == 32'd972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	362   :   assert (rdbk == 32'd3222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	363   :   assert (rdbk == 32'd5209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	364   :   assert (rdbk == 32'd7660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	365   :   assert (rdbk == 32'd11592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	366   :   assert (rdbk == 32'd4965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	367   :   assert (rdbk == 32'd9341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	368   :   assert (rdbk == 32'd526) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	369   :   assert (rdbk == 32'd8664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	370   :   assert (rdbk == 32'd9546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	371   :   assert (rdbk == 32'd1536) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	372   :   assert (rdbk == 32'd3669) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	373   :   assert (rdbk == 32'd11279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	374   :   assert (rdbk == 32'd10845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	375   :   assert (rdbk == 32'd11474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	376   :   assert (rdbk == 32'd10742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	377   :   assert (rdbk == 32'd1391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	378   :   assert (rdbk == 32'd6888) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	379   :   assert (rdbk == 32'd12033) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	380   :   assert (rdbk == 32'd7095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	381   :   assert (rdbk == 32'd8088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	382   :   assert (rdbk == 32'd8931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	383   :   assert (rdbk == 32'd4210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	384   :   assert (rdbk == 32'd7058) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	385   :   assert (rdbk == 32'd3337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	386   :   assert (rdbk == 32'd8259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	387   :   assert (rdbk == 32'd10161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	388   :   assert (rdbk == 32'd12033) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	389   :   assert (rdbk == 32'd6403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	390   :   assert (rdbk == 32'd395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	391   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	392   :   assert (rdbk == 32'd4704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	393   :   assert (rdbk == 32'd976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	394   :   assert (rdbk == 32'd4295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	395   :   assert (rdbk == 32'd1130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	396   :   assert (rdbk == 32'd3146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	397   :   assert (rdbk == 32'd12118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	398   :   assert (rdbk == 32'd7457) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	399   :   assert (rdbk == 32'd12247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	400   :   assert (rdbk == 32'd11727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	401   :   assert (rdbk == 32'd606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	402   :   assert (rdbk == 32'd7340) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	403   :   assert (rdbk == 32'd5760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	404   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	405   :   assert (rdbk == 32'd3991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	406   :   assert (rdbk == 32'd5890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	407   :   assert (rdbk == 32'd3864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	408   :   assert (rdbk == 32'd8942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	409   :   assert (rdbk == 32'd4167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	410   :   assert (rdbk == 32'd10354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	411   :   assert (rdbk == 32'd8794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	412   :   assert (rdbk == 32'd10467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	413   :   assert (rdbk == 32'd1009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	414   :   assert (rdbk == 32'd2762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	415   :   assert (rdbk == 32'd7702) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	416   :   assert (rdbk == 32'd4856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	417   :   assert (rdbk == 32'd1494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	418   :   assert (rdbk == 32'd2156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	419   :   assert (rdbk == 32'd4415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	420   :   assert (rdbk == 32'd6174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	421   :   assert (rdbk == 32'd7215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	422   :   assert (rdbk == 32'd10760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	423   :   assert (rdbk == 32'd10931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	424   :   assert (rdbk == 32'd7300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	425   :   assert (rdbk == 32'd3504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	426   :   assert (rdbk == 32'd4992) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	427   :   assert (rdbk == 32'd10211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	428   :   assert (rdbk == 32'd12172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	429   :   assert (rdbk == 32'd7585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	430   :   assert (rdbk == 32'd4452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	431   :   assert (rdbk == 32'd4010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	432   :   assert (rdbk == 32'd11778) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	433   :   assert (rdbk == 32'd2935) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	434   :   assert (rdbk == 32'd2829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	435   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	436   :   assert (rdbk == 32'd1164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	437   :   assert (rdbk == 32'd5213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	438   :   assert (rdbk == 32'd11522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	439   :   assert (rdbk == 32'd4509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	440   :   assert (rdbk == 32'd10678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	441   :   assert (rdbk == 32'd7847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	442   :   assert (rdbk == 32'd7948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	443   :   assert (rdbk == 32'd5350) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	444   :   assert (rdbk == 32'd1710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	445   :   assert (rdbk == 32'd3253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	446   :   assert (rdbk == 32'd3120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	447   :   assert (rdbk == 32'd1995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	448   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	449   :   assert (rdbk == 32'd3883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	450   :   assert (rdbk == 32'd9425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	451   :   assert (rdbk == 32'd7414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	452   :   assert (rdbk == 32'd803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	453   :   assert (rdbk == 32'd7655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	454   :   assert (rdbk == 32'd10501) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	455   :   assert (rdbk == 32'd6805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	456   :   assert (rdbk == 32'd7214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	457   :   assert (rdbk == 32'd8275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	458   :   assert (rdbk == 32'd1856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	459   :   assert (rdbk == 32'd5480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	460   :   assert (rdbk == 32'd1282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	461   :   assert (rdbk == 32'd9736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	462   :   assert (rdbk == 32'd2185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	463   :   assert (rdbk == 32'd2315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	464   :   assert (rdbk == 32'd2226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	465   :   assert (rdbk == 32'd11611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	466   :   assert (rdbk == 32'd9221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	467   :   assert (rdbk == 32'd10590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	468   :   assert (rdbk == 32'd7730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	469   :   assert (rdbk == 32'd5299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	470   :   assert (rdbk == 32'd6630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	471   :   assert (rdbk == 32'd2380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	472   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	473   :   assert (rdbk == 32'd5278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	474   :   assert (rdbk == 32'd470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	475   :   assert (rdbk == 32'd4668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	476   :   assert (rdbk == 32'd3233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	477   :   assert (rdbk == 32'd1815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	478   :   assert (rdbk == 32'd10840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	479   :   assert (rdbk == 32'd11522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	480   :   assert (rdbk == 32'd3421) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	481   :   assert (rdbk == 32'd5631) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	482   :   assert (rdbk == 32'd11939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	483   :   assert (rdbk == 32'd10708) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	484   :   assert (rdbk == 32'd4709) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	485   :   assert (rdbk == 32'd5447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	486   :   assert (rdbk == 32'd3229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	487   :   assert (rdbk == 32'd8382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	488   :   assert (rdbk == 32'd3826) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	489   :   assert (rdbk == 32'd7791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	490   :   assert (rdbk == 32'd3597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	491   :   assert (rdbk == 32'd8338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	492   :   assert (rdbk == 32'd10040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	493   :   assert (rdbk == 32'd1617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	494   :   assert (rdbk == 32'd1191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	495   :   assert (rdbk == 32'd3678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	496   :   assert (rdbk == 32'd7752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	497   :   assert (rdbk == 32'd4197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	498   :   assert (rdbk == 32'd3100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	499   :   assert (rdbk == 32'd8216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	500   :   assert (rdbk == 32'd7443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	501   :   assert (rdbk == 32'd6488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	502   :   assert (rdbk == 32'd973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	503   :   assert (rdbk == 32'd11347) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	504   :   assert (rdbk == 32'd8865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	505   :   assert (rdbk == 32'd9789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	506   :   assert (rdbk == 32'd1219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	507   :   assert (rdbk == 32'd8020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	508   :   assert (rdbk == 32'd9646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	509   :   assert (rdbk == 32'd9554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	510   :   assert (rdbk == 32'd9786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	511   :   assert (rdbk == 32'd4045) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
    endcase
end


