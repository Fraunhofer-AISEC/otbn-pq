// Copyright Copyright Fraunhofer Institute for Applied and Integrated Security (AISEC).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

$fwrite(f,"----------------------------------------------------------------\n");   
$fwrite(f,"-- PQ-NTT-Indirect (Falcon-1024)\n");
$fwrite(f,"----------------------------------------------------------------\n");   
     
// Write IMEM from File
write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq_ntt_indirect_falcon-1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- IMEM\n");
// Read IMEM  
for (int i=0 ; i<129 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end     

 // Write DMEM from File
write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq_ntt_indirect_falcon-1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

$fwrite(f,"-- DMEM\n");
// Read DMEM  
for (int i=0 ; i<16 ; i++) begin 
    //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
end   
	   
$fwrite(f,"----------------------------------------------------------------\n");   

// Set Instruction Counter to zero (optional)
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );

// Start Programm in IMEM
write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(CmdExecute), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
cc_start = cc;
// Poll on Status Register until Programm is finished
rdbk = '1;
while (rdbk != '0) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
end 

// Measure CC
cc_stop = cc; 
cc_count_falcon1024_indirect = cc_stop - cc_start;        
       
// Read DMEM  
for (int i=0 ; i<1024 ; i++) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+192), .tl_o(tl_o), .tl_i(tl_i_d) );
    
    case(i)
	0   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1   :   assert (rdbk == 32'd969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2   :   assert (rdbk == 32'd5660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3   :   assert (rdbk == 32'd6117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4   :   assert (rdbk == 32'd7575) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	5   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	6   :   assert (rdbk == 32'd11873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	7   :   assert (rdbk == 32'd9428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	8   :   assert (rdbk == 32'd5469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	9   :   assert (rdbk == 32'd5449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	10   :   assert (rdbk == 32'd4522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	11   :   assert (rdbk == 32'd11336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	12   :   assert (rdbk == 32'd1799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	13   :   assert (rdbk == 32'd9101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	14   :   assert (rdbk == 32'd2447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	15   :   assert (rdbk == 32'd2339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	16   :   assert (rdbk == 32'd9415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	17   :   assert (rdbk == 32'd10497) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	18   :   assert (rdbk == 32'd8616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	19   :   assert (rdbk == 32'd11953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	20   :   assert (rdbk == 32'd6800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	21   :   assert (rdbk == 32'd829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	22   :   assert (rdbk == 32'd4677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	23   :   assert (rdbk == 32'd1986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	24   :   assert (rdbk == 32'd4074) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	25   :   assert (rdbk == 32'd2218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	26   :   assert (rdbk == 32'd12162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	27   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	28   :   assert (rdbk == 32'd4464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	29   :   assert (rdbk == 32'd1532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	30   :   assert (rdbk == 32'd2854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	31   :   assert (rdbk == 32'd1578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	32   :   assert (rdbk == 32'd603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	33   :   assert (rdbk == 32'd8964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	34   :   assert (rdbk == 32'd4048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	35   :   assert (rdbk == 32'd5257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	36   :   assert (rdbk == 32'd5925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	37   :   assert (rdbk == 32'd1202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	38   :   assert (rdbk == 32'd5989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	39   :   assert (rdbk == 32'd7571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	40   :   assert (rdbk == 32'd10995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	41   :   assert (rdbk == 32'd2118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	42   :   assert (rdbk == 32'd7621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	43   :   assert (rdbk == 32'd7308) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	44   :   assert (rdbk == 32'd5468) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	45   :   assert (rdbk == 32'd3681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	46   :   assert (rdbk == 32'd3495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	47   :   assert (rdbk == 32'd4090) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	48   :   assert (rdbk == 32'd4201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	49   :   assert (rdbk == 32'd1912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	50   :   assert (rdbk == 32'd11696) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	51   :   assert (rdbk == 32'd8473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	52   :   assert (rdbk == 32'd6720) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	53   :   assert (rdbk == 32'd5259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	54   :   assert (rdbk == 32'd4886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	55   :   assert (rdbk == 32'd10765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	56   :   assert (rdbk == 32'd9283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	57   :   assert (rdbk == 32'd8861) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	58   :   assert (rdbk == 32'd5835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	59   :   assert (rdbk == 32'd3145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	60   :   assert (rdbk == 32'd9065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	61   :   assert (rdbk == 32'd4485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	62   :   assert (rdbk == 32'd7885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	63   :   assert (rdbk == 32'd1456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	64   :   assert (rdbk == 32'd7369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	65   :   assert (rdbk == 32'd409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	66   :   assert (rdbk == 32'd5525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	67   :   assert (rdbk == 32'd2164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	68   :   assert (rdbk == 32'd8590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	69   :   assert (rdbk == 32'd5722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	70   :   assert (rdbk == 32'd3800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	71   :   assert (rdbk == 32'd10000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	72   :   assert (rdbk == 32'd7335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	73   :   assert (rdbk == 32'd2802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	74   :   assert (rdbk == 32'd6125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	75   :   assert (rdbk == 32'd2837) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	76   :   assert (rdbk == 32'd4174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	77   :   assert (rdbk == 32'd4685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	78   :   assert (rdbk == 32'd10259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	79   :   assert (rdbk == 32'd1444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	80   :   assert (rdbk == 32'd546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	81   :   assert (rdbk == 32'd3785) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	82   :   assert (rdbk == 32'd819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	83   :   assert (rdbk == 32'd8037) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	84   :   assert (rdbk == 32'd4567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	85   :   assert (rdbk == 32'd4412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	86   :   assert (rdbk == 32'd1919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	87   :   assert (rdbk == 32'd4691) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	88   :   assert (rdbk == 32'd7804) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	89   :   assert (rdbk == 32'd12106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	90   :   assert (rdbk == 32'd1247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	91   :   assert (rdbk == 32'd2156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	92   :   assert (rdbk == 32'd12180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	93   :   assert (rdbk == 32'd8684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	94   :   assert (rdbk == 32'd5624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	95   :   assert (rdbk == 32'd3071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	96   :   assert (rdbk == 32'd5362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	97   :   assert (rdbk == 32'd4263) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	98   :   assert (rdbk == 32'd11224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	99   :   assert (rdbk == 32'd10223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	100   :   assert (rdbk == 32'd11022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	101   :   assert (rdbk == 32'd3029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	102   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	103   :   assert (rdbk == 32'd9641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	104   :   assert (rdbk == 32'd9815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	105   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	106   :   assert (rdbk == 32'd4010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	107   :   assert (rdbk == 32'd8969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	108   :   assert (rdbk == 32'd7796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	109   :   assert (rdbk == 32'd8428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	110   :   assert (rdbk == 32'd11729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	111   :   assert (rdbk == 32'd2789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	112   :   assert (rdbk == 32'd3569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	113   :   assert (rdbk == 32'd9429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	114   :   assert (rdbk == 32'd11112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	115   :   assert (rdbk == 32'd10591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	116   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	117   :   assert (rdbk == 32'd6909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	118   :   assert (rdbk == 32'd10816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	119   :   assert (rdbk == 32'd768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	120   :   assert (rdbk == 32'd11534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	121   :   assert (rdbk == 32'd8143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	122   :   assert (rdbk == 32'd892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	123   :   assert (rdbk == 32'd6879) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	124   :   assert (rdbk == 32'd11849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	125   :   assert (rdbk == 32'd3624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	126   :   assert (rdbk == 32'd11977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	127   :   assert (rdbk == 32'd5572) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	128   :   assert (rdbk == 32'd4337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	129   :   assert (rdbk == 32'd10647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	130   :   assert (rdbk == 32'd4676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	131   :   assert (rdbk == 32'd8126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	132   :   assert (rdbk == 32'd5777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	133   :   assert (rdbk == 32'd3496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	134   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	135   :   assert (rdbk == 32'd405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	136   :   assert (rdbk == 32'd6375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	137   :   assert (rdbk == 32'd1599) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	138   :   assert (rdbk == 32'd2625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	139   :   assert (rdbk == 32'd6154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	140   :   assert (rdbk == 32'd2253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	141   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	142   :   assert (rdbk == 32'd931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	143   :   assert (rdbk == 32'd11330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	144   :   assert (rdbk == 32'd1184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	145   :   assert (rdbk == 32'd2936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	146   :   assert (rdbk == 32'd1563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	147   :   assert (rdbk == 32'd11379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	148   :   assert (rdbk == 32'd8515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	149   :   assert (rdbk == 32'd8066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	150   :   assert (rdbk == 32'd9978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	151   :   assert (rdbk == 32'd9988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	152   :   assert (rdbk == 32'd10979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	153   :   assert (rdbk == 32'd5467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	154   :   assert (rdbk == 32'd1401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	155   :   assert (rdbk == 32'd6246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	156   :   assert (rdbk == 32'd12144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	157   :   assert (rdbk == 32'd11241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	158   :   assert (rdbk == 32'd3840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	159   :   assert (rdbk == 32'd3627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	160   :   assert (rdbk == 32'd2936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	161   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	162   :   assert (rdbk == 32'd948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	163   :   assert (rdbk == 32'd7804) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	164   :   assert (rdbk == 32'd10522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	165   :   assert (rdbk == 32'd2546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	166   :   assert (rdbk == 32'd687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	167   :   assert (rdbk == 32'd532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	168   :   assert (rdbk == 32'd8222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	169   :   assert (rdbk == 32'd10937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	170   :   assert (rdbk == 32'd545) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	171   :   assert (rdbk == 32'd6775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	172   :   assert (rdbk == 32'd12003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	173   :   assert (rdbk == 32'd336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	174   :   assert (rdbk == 32'd9381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	175   :   assert (rdbk == 32'd6279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	176   :   assert (rdbk == 32'd4028) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	177   :   assert (rdbk == 32'd8884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	178   :   assert (rdbk == 32'd11513) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	179   :   assert (rdbk == 32'd3383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	180   :   assert (rdbk == 32'd3204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	181   :   assert (rdbk == 32'd4385) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	182   :   assert (rdbk == 32'd1425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	183   :   assert (rdbk == 32'd6394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	184   :   assert (rdbk == 32'd8439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	185   :   assert (rdbk == 32'd5251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	186   :   assert (rdbk == 32'd11056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	187   :   assert (rdbk == 32'd5140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	188   :   assert (rdbk == 32'd4397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	189   :   assert (rdbk == 32'd6355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	190   :   assert (rdbk == 32'd8557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	191   :   assert (rdbk == 32'd12271) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	192   :   assert (rdbk == 32'd12081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	193   :   assert (rdbk == 32'd5791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	194   :   assert (rdbk == 32'd2115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	195   :   assert (rdbk == 32'd10144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	196   :   assert (rdbk == 32'd9144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	197   :   assert (rdbk == 32'd5406) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	198   :   assert (rdbk == 32'd6557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	199   :   assert (rdbk == 32'd1557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	200   :   assert (rdbk == 32'd2169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	201   :   assert (rdbk == 32'd5148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	202   :   assert (rdbk == 32'd11654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	203   :   assert (rdbk == 32'd6500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	204   :   assert (rdbk == 32'd7105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	205   :   assert (rdbk == 32'd3905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	206   :   assert (rdbk == 32'd11692) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	207   :   assert (rdbk == 32'd1038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	208   :   assert (rdbk == 32'd5949) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	209   :   assert (rdbk == 32'd10896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	210   :   assert (rdbk == 32'd9340) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	211   :   assert (rdbk == 32'd1946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	212   :   assert (rdbk == 32'd8715) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	213   :   assert (rdbk == 32'd11530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	214   :   assert (rdbk == 32'd8030) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	215   :   assert (rdbk == 32'd2904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	216   :   assert (rdbk == 32'd9384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	217   :   assert (rdbk == 32'd8968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	218   :   assert (rdbk == 32'd5281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	219   :   assert (rdbk == 32'd2884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	220   :   assert (rdbk == 32'd9286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	221   :   assert (rdbk == 32'd6884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	222   :   assert (rdbk == 32'd1179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	223   :   assert (rdbk == 32'd1444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	224   :   assert (rdbk == 32'd4934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	225   :   assert (rdbk == 32'd3832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	226   :   assert (rdbk == 32'd11104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	227   :   assert (rdbk == 32'd4933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	228   :   assert (rdbk == 32'd6958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	229   :   assert (rdbk == 32'd8752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	230   :   assert (rdbk == 32'd9820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	231   :   assert (rdbk == 32'd719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	232   :   assert (rdbk == 32'd9763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	233   :   assert (rdbk == 32'd6140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	234   :   assert (rdbk == 32'd848) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	235   :   assert (rdbk == 32'd836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	236   :   assert (rdbk == 32'd11737) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	237   :   assert (rdbk == 32'd8942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	238   :   assert (rdbk == 32'd1793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	239   :   assert (rdbk == 32'd6901) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	240   :   assert (rdbk == 32'd6989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	241   :   assert (rdbk == 32'd11926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	242   :   assert (rdbk == 32'd6004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	243   :   assert (rdbk == 32'd1571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	244   :   assert (rdbk == 32'd7780) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	245   :   assert (rdbk == 32'd9774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	246   :   assert (rdbk == 32'd412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	247   :   assert (rdbk == 32'd3001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	248   :   assert (rdbk == 32'd3558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	249   :   assert (rdbk == 32'd579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	250   :   assert (rdbk == 32'd4020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	251   :   assert (rdbk == 32'd7384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	252   :   assert (rdbk == 32'd6341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	253   :   assert (rdbk == 32'd11712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	254   :   assert (rdbk == 32'd9904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	255   :   assert (rdbk == 32'd4976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	256   :   assert (rdbk == 32'd547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	257   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	258   :   assert (rdbk == 32'd6409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	259   :   assert (rdbk == 32'd10437) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	260   :   assert (rdbk == 32'd11494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	261   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	262   :   assert (rdbk == 32'd9789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	263   :   assert (rdbk == 32'd2325) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	264   :   assert (rdbk == 32'd1314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	265   :   assert (rdbk == 32'd2516) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	266   :   assert (rdbk == 32'd6846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	267   :   assert (rdbk == 32'd8870) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	268   :   assert (rdbk == 32'd11616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	269   :   assert (rdbk == 32'd10635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	270   :   assert (rdbk == 32'd5621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	271   :   assert (rdbk == 32'd9665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	272   :   assert (rdbk == 32'd3189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	273   :   assert (rdbk == 32'd4624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	274   :   assert (rdbk == 32'd718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	275   :   assert (rdbk == 32'd9494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	276   :   assert (rdbk == 32'd12124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	277   :   assert (rdbk == 32'd3016) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	278   :   assert (rdbk == 32'd7819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	279   :   assert (rdbk == 32'd11466) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	280   :   assert (rdbk == 32'd825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	281   :   assert (rdbk == 32'd11349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	282   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	283   :   assert (rdbk == 32'd1739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	284   :   assert (rdbk == 32'd11141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	285   :   assert (rdbk == 32'd8021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	286   :   assert (rdbk == 32'd7381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	287   :   assert (rdbk == 32'd3759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	288   :   assert (rdbk == 32'd11968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	289   :   assert (rdbk == 32'd9622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	290   :   assert (rdbk == 32'd10046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	291   :   assert (rdbk == 32'd9282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	292   :   assert (rdbk == 32'd10881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	293   :   assert (rdbk == 32'd1533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	294   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	295   :   assert (rdbk == 32'd8763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	296   :   assert (rdbk == 32'd8758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	297   :   assert (rdbk == 32'd2219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	298   :   assert (rdbk == 32'd11566) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	299   :   assert (rdbk == 32'd9225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	300   :   assert (rdbk == 32'd899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	301   :   assert (rdbk == 32'd10687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	302   :   assert (rdbk == 32'd9761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	303   :   assert (rdbk == 32'd8476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	304   :   assert (rdbk == 32'd782) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	305   :   assert (rdbk == 32'd8964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	306   :   assert (rdbk == 32'd3707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	307   :   assert (rdbk == 32'd4916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	308   :   assert (rdbk == 32'd1344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	309   :   assert (rdbk == 32'd10994) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	310   :   assert (rdbk == 32'd12098) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	311   :   assert (rdbk == 32'd9963) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	312   :   assert (rdbk == 32'd1833) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	313   :   assert (rdbk == 32'd2509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	314   :   assert (rdbk == 32'd7758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	315   :   assert (rdbk == 32'd1720) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	316   :   assert (rdbk == 32'd2362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	317   :   assert (rdbk == 32'd4802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	318   :   assert (rdbk == 32'd9733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	319   :   assert (rdbk == 32'd3989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	320   :   assert (rdbk == 32'd8666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	321   :   assert (rdbk == 32'd9946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	322   :   assert (rdbk == 32'd1489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	323   :   assert (rdbk == 32'd3299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	324   :   assert (rdbk == 32'd5017) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	325   :   assert (rdbk == 32'd3117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	326   :   assert (rdbk == 32'd3431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	327   :   assert (rdbk == 32'd5550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	328   :   assert (rdbk == 32'd1755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	329   :   assert (rdbk == 32'd9313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	330   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	331   :   assert (rdbk == 32'd1581) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	332   :   assert (rdbk == 32'd8624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	333   :   assert (rdbk == 32'd2355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	334   :   assert (rdbk == 32'd772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	335   :   assert (rdbk == 32'd9783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	336   :   assert (rdbk == 32'd10114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	337   :   assert (rdbk == 32'd5276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	338   :   assert (rdbk == 32'd786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	339   :   assert (rdbk == 32'd10628) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	340   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	341   :   assert (rdbk == 32'd3420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	342   :   assert (rdbk == 32'd4101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	343   :   assert (rdbk == 32'd10850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	344   :   assert (rdbk == 32'd5560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	345   :   assert (rdbk == 32'd2035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	346   :   assert (rdbk == 32'd9111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	347   :   assert (rdbk == 32'd1100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	348   :   assert (rdbk == 32'd4239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	349   :   assert (rdbk == 32'd7282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	350   :   assert (rdbk == 32'd2398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	351   :   assert (rdbk == 32'd2881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	352   :   assert (rdbk == 32'd10485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	353   :   assert (rdbk == 32'd3639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	354   :   assert (rdbk == 32'd11057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	355   :   assert (rdbk == 32'd10188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	356   :   assert (rdbk == 32'd1531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	357   :   assert (rdbk == 32'd9694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	358   :   assert (rdbk == 32'd11605) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	359   :   assert (rdbk == 32'd2151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	360   :   assert (rdbk == 32'd9062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	361   :   assert (rdbk == 32'd8570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	362   :   assert (rdbk == 32'd9294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	363   :   assert (rdbk == 32'd1307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	364   :   assert (rdbk == 32'd2452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	365   :   assert (rdbk == 32'd11202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	366   :   assert (rdbk == 32'd2618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	367   :   assert (rdbk == 32'd1703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	368   :   assert (rdbk == 32'd7979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	369   :   assert (rdbk == 32'd6564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	370   :   assert (rdbk == 32'd5309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	371   :   assert (rdbk == 32'd4351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	372   :   assert (rdbk == 32'd5578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	373   :   assert (rdbk == 32'd11815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	374   :   assert (rdbk == 32'd4805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	375   :   assert (rdbk == 32'd11952) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	376   :   assert (rdbk == 32'd6307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	377   :   assert (rdbk == 32'd11363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	378   :   assert (rdbk == 32'd8394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	379   :   assert (rdbk == 32'd11307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	380   :   assert (rdbk == 32'd5817) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	381   :   assert (rdbk == 32'd2972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	382   :   assert (rdbk == 32'd10746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	383   :   assert (rdbk == 32'd3724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	384   :   assert (rdbk == 32'd11492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	385   :   assert (rdbk == 32'd10863) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	386   :   assert (rdbk == 32'd965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	387   :   assert (rdbk == 32'd5598) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	388   :   assert (rdbk == 32'd3117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	389   :   assert (rdbk == 32'd5874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	390   :   assert (rdbk == 32'd7251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	391   :   assert (rdbk == 32'd3264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	392   :   assert (rdbk == 32'd619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	393   :   assert (rdbk == 32'd6646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	394   :   assert (rdbk == 32'd1669) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	395   :   assert (rdbk == 32'd10024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	396   :   assert (rdbk == 32'd11174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	397   :   assert (rdbk == 32'd8099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	398   :   assert (rdbk == 32'd6001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	399   :   assert (rdbk == 32'd8416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	400   :   assert (rdbk == 32'd6640) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	401   :   assert (rdbk == 32'd10945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	402   :   assert (rdbk == 32'd6446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	403   :   assert (rdbk == 32'd10580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	404   :   assert (rdbk == 32'd4182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	405   :   assert (rdbk == 32'd8414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	406   :   assert (rdbk == 32'd6024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	407   :   assert (rdbk == 32'd3368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	408   :   assert (rdbk == 32'd10066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	409   :   assert (rdbk == 32'd8153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	410   :   assert (rdbk == 32'd634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	411   :   assert (rdbk == 32'd6099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	412   :   assert (rdbk == 32'd1288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	413   :   assert (rdbk == 32'd4330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	414   :   assert (rdbk == 32'd4394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	415   :   assert (rdbk == 32'd1483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	416   :   assert (rdbk == 32'd8290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	417   :   assert (rdbk == 32'd865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	418   :   assert (rdbk == 32'd8113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	419   :   assert (rdbk == 32'd965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	420   :   assert (rdbk == 32'd12022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	421   :   assert (rdbk == 32'd10529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	422   :   assert (rdbk == 32'd5638) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	423   :   assert (rdbk == 32'd7321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	424   :   assert (rdbk == 32'd2972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	425   :   assert (rdbk == 32'd3571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	426   :   assert (rdbk == 32'd3039) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	427   :   assert (rdbk == 32'd6356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	428   :   assert (rdbk == 32'd11008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	429   :   assert (rdbk == 32'd6124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	430   :   assert (rdbk == 32'd6452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	431   :   assert (rdbk == 32'd6926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	432   :   assert (rdbk == 32'd8061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	433   :   assert (rdbk == 32'd9565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	434   :   assert (rdbk == 32'd9356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	435   :   assert (rdbk == 32'd3929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	436   :   assert (rdbk == 32'd3318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	437   :   assert (rdbk == 32'd7265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	438   :   assert (rdbk == 32'd4468) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	439   :   assert (rdbk == 32'd9710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	440   :   assert (rdbk == 32'd4803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	441   :   assert (rdbk == 32'd4770) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	442   :   assert (rdbk == 32'd6579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	443   :   assert (rdbk == 32'd5071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	444   :   assert (rdbk == 32'd2982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	445   :   assert (rdbk == 32'd1497) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	446   :   assert (rdbk == 32'd10113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	447   :   assert (rdbk == 32'd4482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	448   :   assert (rdbk == 32'd9682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	449   :   assert (rdbk == 32'd11039) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	450   :   assert (rdbk == 32'd7354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	451   :   assert (rdbk == 32'd8436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	452   :   assert (rdbk == 32'd5665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	453   :   assert (rdbk == 32'd2869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	454   :   assert (rdbk == 32'd7998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	455   :   assert (rdbk == 32'd5718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	456   :   assert (rdbk == 32'd9467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	457   :   assert (rdbk == 32'd3749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	458   :   assert (rdbk == 32'd4956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	459   :   assert (rdbk == 32'd8447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	460   :   assert (rdbk == 32'd10496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	461   :   assert (rdbk == 32'd11803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	462   :   assert (rdbk == 32'd10627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	463   :   assert (rdbk == 32'd10102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	464   :   assert (rdbk == 32'd7682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	465   :   assert (rdbk == 32'd1277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	466   :   assert (rdbk == 32'd4255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	467   :   assert (rdbk == 32'd11229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	468   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	469   :   assert (rdbk == 32'd7627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	470   :   assert (rdbk == 32'd6936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	471   :   assert (rdbk == 32'd3027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	472   :   assert (rdbk == 32'd2515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	473   :   assert (rdbk == 32'd2339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	474   :   assert (rdbk == 32'd7313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	475   :   assert (rdbk == 32'd2851) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	476   :   assert (rdbk == 32'd5346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	477   :   assert (rdbk == 32'd1481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	478   :   assert (rdbk == 32'd8854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	479   :   assert (rdbk == 32'd7341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	480   :   assert (rdbk == 32'd10075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	481   :   assert (rdbk == 32'd3191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	482   :   assert (rdbk == 32'd4110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	483   :   assert (rdbk == 32'd7843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	484   :   assert (rdbk == 32'd10609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	485   :   assert (rdbk == 32'd10343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	486   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	487   :   assert (rdbk == 32'd4885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	488   :   assert (rdbk == 32'd3771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	489   :   assert (rdbk == 32'd11524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	490   :   assert (rdbk == 32'd8472) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	491   :   assert (rdbk == 32'd2623) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	492   :   assert (rdbk == 32'd10040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	493   :   assert (rdbk == 32'd7927) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	494   :   assert (rdbk == 32'd7400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	495   :   assert (rdbk == 32'd660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	496   :   assert (rdbk == 32'd1585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	497   :   assert (rdbk == 32'd11891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	498   :   assert (rdbk == 32'd9882) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	499   :   assert (rdbk == 32'd724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	500   :   assert (rdbk == 32'd4854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	501   :   assert (rdbk == 32'd3823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	502   :   assert (rdbk == 32'd4109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	503   :   assert (rdbk == 32'd3192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	504   :   assert (rdbk == 32'd5359) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	505   :   assert (rdbk == 32'd8327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	506   :   assert (rdbk == 32'd4241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	507   :   assert (rdbk == 32'd1990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	508   :   assert (rdbk == 32'd7253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	509   :   assert (rdbk == 32'd274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	510   :   assert (rdbk == 32'd2010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	511   :   assert (rdbk == 32'd2346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	512   :   assert (rdbk == 32'd4566) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	513   :   assert (rdbk == 32'd9384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	514   :   assert (rdbk == 32'd997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	515   :   assert (rdbk == 32'd7425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	516   :   assert (rdbk == 32'd2619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	517   :   assert (rdbk == 32'd7567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	518   :   assert (rdbk == 32'd7740) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	519   :   assert (rdbk == 32'd1981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	520   :   assert (rdbk == 32'd2357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	521   :   assert (rdbk == 32'd7122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	522   :   assert (rdbk == 32'd9314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	523   :   assert (rdbk == 32'd7314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	524   :   assert (rdbk == 32'd9945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	525   :   assert (rdbk == 32'd4561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	526   :   assert (rdbk == 32'd6611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	527   :   assert (rdbk == 32'd5827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	528   :   assert (rdbk == 32'd4027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	529   :   assert (rdbk == 32'd10647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	530   :   assert (rdbk == 32'd5377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	531   :   assert (rdbk == 32'd4841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	532   :   assert (rdbk == 32'd12169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	533   :   assert (rdbk == 32'd9494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	534   :   assert (rdbk == 32'd8503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	535   :   assert (rdbk == 32'd3571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	536   :   assert (rdbk == 32'd3579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	537   :   assert (rdbk == 32'd1794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	538   :   assert (rdbk == 32'd5911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	539   :   assert (rdbk == 32'd3317) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	540   :   assert (rdbk == 32'd1971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	541   :   assert (rdbk == 32'd5904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	542   :   assert (rdbk == 32'd6239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	543   :   assert (rdbk == 32'd2867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	544   :   assert (rdbk == 32'd5239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	545   :   assert (rdbk == 32'd4982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	546   :   assert (rdbk == 32'd267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	547   :   assert (rdbk == 32'd5836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	548   :   assert (rdbk == 32'd10102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	549   :   assert (rdbk == 32'd7324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	550   :   assert (rdbk == 32'd7778) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	551   :   assert (rdbk == 32'd3086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	552   :   assert (rdbk == 32'd6484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	553   :   assert (rdbk == 32'd6379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	554   :   assert (rdbk == 32'd4448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	555   :   assert (rdbk == 32'd3228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	556   :   assert (rdbk == 32'd9764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	557   :   assert (rdbk == 32'd7514) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	558   :   assert (rdbk == 32'd931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	559   :   assert (rdbk == 32'd8067) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	560   :   assert (rdbk == 32'd7876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	561   :   assert (rdbk == 32'd4961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	562   :   assert (rdbk == 32'd1621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	563   :   assert (rdbk == 32'd1743) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	564   :   assert (rdbk == 32'd1743) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	565   :   assert (rdbk == 32'd11298) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	566   :   assert (rdbk == 32'd2953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	567   :   assert (rdbk == 32'd2871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	568   :   assert (rdbk == 32'd677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	569   :   assert (rdbk == 32'd11476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	570   :   assert (rdbk == 32'd6086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	571   :   assert (rdbk == 32'd8758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	572   :   assert (rdbk == 32'd7723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	573   :   assert (rdbk == 32'd1461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	574   :   assert (rdbk == 32'd6739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	575   :   assert (rdbk == 32'd11664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	576   :   assert (rdbk == 32'd9763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	577   :   assert (rdbk == 32'd8570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	578   :   assert (rdbk == 32'd373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	579   :   assert (rdbk == 32'd5812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	580   :   assert (rdbk == 32'd5462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	581   :   assert (rdbk == 32'd746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	582   :   assert (rdbk == 32'd6093) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	583   :   assert (rdbk == 32'd1665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	584   :   assert (rdbk == 32'd5289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	585   :   assert (rdbk == 32'd3846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	586   :   assert (rdbk == 32'd6630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	587   :   assert (rdbk == 32'd5182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	588   :   assert (rdbk == 32'd3897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	589   :   assert (rdbk == 32'd7075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	590   :   assert (rdbk == 32'd8970) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	591   :   assert (rdbk == 32'd10147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	592   :   assert (rdbk == 32'd5481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	593   :   assert (rdbk == 32'd7667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	594   :   assert (rdbk == 32'd11083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	595   :   assert (rdbk == 32'd3966) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	596   :   assert (rdbk == 32'd5283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	597   :   assert (rdbk == 32'd6106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	598   :   assert (rdbk == 32'd4232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	599   :   assert (rdbk == 32'd3084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	600   :   assert (rdbk == 32'd4998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	601   :   assert (rdbk == 32'd1314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	602   :   assert (rdbk == 32'd3636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	603   :   assert (rdbk == 32'd11856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	604   :   assert (rdbk == 32'd8397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	605   :   assert (rdbk == 32'd7463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	606   :   assert (rdbk == 32'd4532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	607   :   assert (rdbk == 32'd5219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	608   :   assert (rdbk == 32'd6511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	609   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	610   :   assert (rdbk == 32'd7849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	611   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	612   :   assert (rdbk == 32'd8807) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	613   :   assert (rdbk == 32'd1984) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	614   :   assert (rdbk == 32'd8233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	615   :   assert (rdbk == 32'd3761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	616   :   assert (rdbk == 32'd1024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	617   :   assert (rdbk == 32'd8529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	618   :   assert (rdbk == 32'd1259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	619   :   assert (rdbk == 32'd9393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	620   :   assert (rdbk == 32'd6759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	621   :   assert (rdbk == 32'd1568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	622   :   assert (rdbk == 32'd5187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	623   :   assert (rdbk == 32'd10634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	624   :   assert (rdbk == 32'd9245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	625   :   assert (rdbk == 32'd3215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	626   :   assert (rdbk == 32'd11521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	627   :   assert (rdbk == 32'd9348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	628   :   assert (rdbk == 32'd8820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	629   :   assert (rdbk == 32'd7716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	630   :   assert (rdbk == 32'd8371) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	631   :   assert (rdbk == 32'd7655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	632   :   assert (rdbk == 32'd1914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	633   :   assert (rdbk == 32'd2644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	634   :   assert (rdbk == 32'd4243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	635   :   assert (rdbk == 32'd1638) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	636   :   assert (rdbk == 32'd2354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	637   :   assert (rdbk == 32'd8712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	638   :   assert (rdbk == 32'd300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	639   :   assert (rdbk == 32'd8305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	640   :   assert (rdbk == 32'd3089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	641   :   assert (rdbk == 32'd8828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	642   :   assert (rdbk == 32'd5856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	643   :   assert (rdbk == 32'd858) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	644   :   assert (rdbk == 32'd4477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	645   :   assert (rdbk == 32'd2567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	646   :   assert (rdbk == 32'd10680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	647   :   assert (rdbk == 32'd2467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	648   :   assert (rdbk == 32'd9065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	649   :   assert (rdbk == 32'd7906) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	650   :   assert (rdbk == 32'd2342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	651   :   assert (rdbk == 32'd7567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	652   :   assert (rdbk == 32'd483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	653   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	654   :   assert (rdbk == 32'd257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	655   :   assert (rdbk == 32'd11499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	656   :   assert (rdbk == 32'd6616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	657   :   assert (rdbk == 32'd2870) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	658   :   assert (rdbk == 32'd12113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	659   :   assert (rdbk == 32'd5554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	660   :   assert (rdbk == 32'd9996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	661   :   assert (rdbk == 32'd9207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	662   :   assert (rdbk == 32'd4630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	663   :   assert (rdbk == 32'd7392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	664   :   assert (rdbk == 32'd4167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	665   :   assert (rdbk == 32'd10276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	666   :   assert (rdbk == 32'd11658) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	667   :   assert (rdbk == 32'd9667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	668   :   assert (rdbk == 32'd5247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	669   :   assert (rdbk == 32'd10030) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	670   :   assert (rdbk == 32'd4814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	671   :   assert (rdbk == 32'd12234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	672   :   assert (rdbk == 32'd6678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	673   :   assert (rdbk == 32'd696) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	674   :   assert (rdbk == 32'd10155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	675   :   assert (rdbk == 32'd2740) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	676   :   assert (rdbk == 32'd2582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	677   :   assert (rdbk == 32'd11793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	678   :   assert (rdbk == 32'd3161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	679   :   assert (rdbk == 32'd3413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	680   :   assert (rdbk == 32'd10981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	681   :   assert (rdbk == 32'd6885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	682   :   assert (rdbk == 32'd11440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	683   :   assert (rdbk == 32'd511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	684   :   assert (rdbk == 32'd3726) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	685   :   assert (rdbk == 32'd3649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	686   :   assert (rdbk == 32'd11686) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	687   :   assert (rdbk == 32'd10147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	688   :   assert (rdbk == 32'd5641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	689   :   assert (rdbk == 32'd12152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	690   :   assert (rdbk == 32'd10550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	691   :   assert (rdbk == 32'd11544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	692   :   assert (rdbk == 32'd8848) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	693   :   assert (rdbk == 32'd381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	694   :   assert (rdbk == 32'd979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	695   :   assert (rdbk == 32'd5847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	696   :   assert (rdbk == 32'd11590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	697   :   assert (rdbk == 32'd7655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	698   :   assert (rdbk == 32'd951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	699   :   assert (rdbk == 32'd8417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	700   :   assert (rdbk == 32'd9096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	701   :   assert (rdbk == 32'd10900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	702   :   assert (rdbk == 32'd8126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	703   :   assert (rdbk == 32'd2962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	704   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	705   :   assert (rdbk == 32'd10767) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	706   :   assert (rdbk == 32'd8559) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	707   :   assert (rdbk == 32'd9181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	708   :   assert (rdbk == 32'd12232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	709   :   assert (rdbk == 32'd11077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	710   :   assert (rdbk == 32'd4563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	711   :   assert (rdbk == 32'd12232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	712   :   assert (rdbk == 32'd275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	713   :   assert (rdbk == 32'd5106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	714   :   assert (rdbk == 32'd1296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	715   :   assert (rdbk == 32'd9180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	716   :   assert (rdbk == 32'd1032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	717   :   assert (rdbk == 32'd11960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	718   :   assert (rdbk == 32'd5312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	719   :   assert (rdbk == 32'd419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	720   :   assert (rdbk == 32'd7311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	721   :   assert (rdbk == 32'd10911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	722   :   assert (rdbk == 32'd11165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	723   :   assert (rdbk == 32'd4435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	724   :   assert (rdbk == 32'd3750) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	725   :   assert (rdbk == 32'd4521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	726   :   assert (rdbk == 32'd11119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	727   :   assert (rdbk == 32'd4012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	728   :   assert (rdbk == 32'd5070) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	729   :   assert (rdbk == 32'd6650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	730   :   assert (rdbk == 32'd10616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	731   :   assert (rdbk == 32'd2061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	732   :   assert (rdbk == 32'd10680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	733   :   assert (rdbk == 32'd6930) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	734   :   assert (rdbk == 32'd7706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	735   :   assert (rdbk == 32'd6985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	736   :   assert (rdbk == 32'd6417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	737   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	738   :   assert (rdbk == 32'd7287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	739   :   assert (rdbk == 32'd10529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	740   :   assert (rdbk == 32'd7219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	741   :   assert (rdbk == 32'd1634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	742   :   assert (rdbk == 32'd5891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	743   :   assert (rdbk == 32'd2208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	744   :   assert (rdbk == 32'd11568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	745   :   assert (rdbk == 32'd6189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	746   :   assert (rdbk == 32'd2119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	747   :   assert (rdbk == 32'd5895) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	748   :   assert (rdbk == 32'd7544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	749   :   assert (rdbk == 32'd991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	750   :   assert (rdbk == 32'd4339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	751   :   assert (rdbk == 32'd3685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	752   :   assert (rdbk == 32'd2121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	753   :   assert (rdbk == 32'd8753) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	754   :   assert (rdbk == 32'd4048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	755   :   assert (rdbk == 32'd6846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	756   :   assert (rdbk == 32'd5681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	757   :   assert (rdbk == 32'd6881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	758   :   assert (rdbk == 32'd9477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	759   :   assert (rdbk == 32'd10942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	760   :   assert (rdbk == 32'd9380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	761   :   assert (rdbk == 32'd273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	762   :   assert (rdbk == 32'd5278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	763   :   assert (rdbk == 32'd3582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	764   :   assert (rdbk == 32'd7958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	765   :   assert (rdbk == 32'd6407) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	766   :   assert (rdbk == 32'd9539) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	767   :   assert (rdbk == 32'd4727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	768   :   assert (rdbk == 32'd919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	769   :   assert (rdbk == 32'd816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	770   :   assert (rdbk == 32'd10272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	771   :   assert (rdbk == 32'd10916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	772   :   assert (rdbk == 32'd1701) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	773   :   assert (rdbk == 32'd4988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	774   :   assert (rdbk == 32'd6354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	775   :   assert (rdbk == 32'd680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	776   :   assert (rdbk == 32'd11504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	777   :   assert (rdbk == 32'd8218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	778   :   assert (rdbk == 32'd11557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	779   :   assert (rdbk == 32'd9012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	780   :   assert (rdbk == 32'd9003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	781   :   assert (rdbk == 32'd10068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	782   :   assert (rdbk == 32'd7205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	783   :   assert (rdbk == 32'd2845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	784   :   assert (rdbk == 32'd8731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	785   :   assert (rdbk == 32'd8122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	786   :   assert (rdbk == 32'd4167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	787   :   assert (rdbk == 32'd6881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	788   :   assert (rdbk == 32'd9430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	789   :   assert (rdbk == 32'd11557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	790   :   assert (rdbk == 32'd9823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	791   :   assert (rdbk == 32'd10649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	792   :   assert (rdbk == 32'd7192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	793   :   assert (rdbk == 32'd2355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	794   :   assert (rdbk == 32'd448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	795   :   assert (rdbk == 32'd3547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	796   :   assert (rdbk == 32'd3095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	797   :   assert (rdbk == 32'd5307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	798   :   assert (rdbk == 32'd3361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	799   :   assert (rdbk == 32'd6225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	800   :   assert (rdbk == 32'd11565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	801   :   assert (rdbk == 32'd7951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	802   :   assert (rdbk == 32'd4476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	803   :   assert (rdbk == 32'd10055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	804   :   assert (rdbk == 32'd4380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	805   :   assert (rdbk == 32'd1212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	806   :   assert (rdbk == 32'd9560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	807   :   assert (rdbk == 32'd6651) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	808   :   assert (rdbk == 32'd3403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	809   :   assert (rdbk == 32'd5777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	810   :   assert (rdbk == 32'd7708) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	811   :   assert (rdbk == 32'd299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	812   :   assert (rdbk == 32'd5364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	813   :   assert (rdbk == 32'd3352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	814   :   assert (rdbk == 32'd9207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	815   :   assert (rdbk == 32'd5304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	816   :   assert (rdbk == 32'd10540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	817   :   assert (rdbk == 32'd10257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	818   :   assert (rdbk == 32'd1768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	819   :   assert (rdbk == 32'd7014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	820   :   assert (rdbk == 32'd1921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	821   :   assert (rdbk == 32'd10607) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	822   :   assert (rdbk == 32'd9384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	823   :   assert (rdbk == 32'd10657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	824   :   assert (rdbk == 32'd10948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	825   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	826   :   assert (rdbk == 32'd5291) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	827   :   assert (rdbk == 32'd7395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	828   :   assert (rdbk == 32'd5916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	829   :   assert (rdbk == 32'd9887) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	830   :   assert (rdbk == 32'd417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	831   :   assert (rdbk == 32'd5760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	832   :   assert (rdbk == 32'd6027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	833   :   assert (rdbk == 32'd1562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	834   :   assert (rdbk == 32'd4114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	835   :   assert (rdbk == 32'd6746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	836   :   assert (rdbk == 32'd9680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	837   :   assert (rdbk == 32'd6129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	838   :   assert (rdbk == 32'd8003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	839   :   assert (rdbk == 32'd5233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	840   :   assert (rdbk == 32'd1495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	841   :   assert (rdbk == 32'd4645) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	842   :   assert (rdbk == 32'd4752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	843   :   assert (rdbk == 32'd11487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	844   :   assert (rdbk == 32'd755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	845   :   assert (rdbk == 32'd8890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	846   :   assert (rdbk == 32'd4126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	847   :   assert (rdbk == 32'd5381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	848   :   assert (rdbk == 32'd4723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	849   :   assert (rdbk == 32'd1837) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	850   :   assert (rdbk == 32'd11599) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	851   :   assert (rdbk == 32'd5527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	852   :   assert (rdbk == 32'd1137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	853   :   assert (rdbk == 32'd11898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	854   :   assert (rdbk == 32'd3503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	855   :   assert (rdbk == 32'd5542) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	856   :   assert (rdbk == 32'd5065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	857   :   assert (rdbk == 32'd2144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	858   :   assert (rdbk == 32'd2351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	859   :   assert (rdbk == 32'd6358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	860   :   assert (rdbk == 32'd11126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	861   :   assert (rdbk == 32'd1681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	862   :   assert (rdbk == 32'd2742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	863   :   assert (rdbk == 32'd5199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	864   :   assert (rdbk == 32'd5720) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	865   :   assert (rdbk == 32'd9439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	866   :   assert (rdbk == 32'd10943) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	867   :   assert (rdbk == 32'd10208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	868   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	869   :   assert (rdbk == 32'd8666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	870   :   assert (rdbk == 32'd11895) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	871   :   assert (rdbk == 32'd1073) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	872   :   assert (rdbk == 32'd1795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	873   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	874   :   assert (rdbk == 32'd8664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	875   :   assert (rdbk == 32'd2892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	876   :   assert (rdbk == 32'd6747) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	877   :   assert (rdbk == 32'd2029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	878   :   assert (rdbk == 32'd6024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	879   :   assert (rdbk == 32'd11867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	880   :   assert (rdbk == 32'd7355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	881   :   assert (rdbk == 32'd5503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	882   :   assert (rdbk == 32'd1441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	883   :   assert (rdbk == 32'd7953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	884   :   assert (rdbk == 32'd6012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	885   :   assert (rdbk == 32'd2726) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	886   :   assert (rdbk == 32'd6583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	887   :   assert (rdbk == 32'd7731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	888   :   assert (rdbk == 32'd3015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	889   :   assert (rdbk == 32'd7420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	890   :   assert (rdbk == 32'd1902) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	891   :   assert (rdbk == 32'd11923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	892   :   assert (rdbk == 32'd10773) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	893   :   assert (rdbk == 32'd10206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	894   :   assert (rdbk == 32'd11656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	895   :   assert (rdbk == 32'd3257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	896   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	897   :   assert (rdbk == 32'd10357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	898   :   assert (rdbk == 32'd268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	899   :   assert (rdbk == 32'd8695) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	900   :   assert (rdbk == 32'd8445) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	901   :   assert (rdbk == 32'd1268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	902   :   assert (rdbk == 32'd11945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	903   :   assert (rdbk == 32'd8144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	904   :   assert (rdbk == 32'd11254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	905   :   assert (rdbk == 32'd10123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	906   :   assert (rdbk == 32'd7628) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	907   :   assert (rdbk == 32'd5082) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	908   :   assert (rdbk == 32'd8264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	909   :   assert (rdbk == 32'd994) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	910   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	911   :   assert (rdbk == 32'd7201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	912   :   assert (rdbk == 32'd6158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	913   :   assert (rdbk == 32'd1825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	914   :   assert (rdbk == 32'd6382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	915   :   assert (rdbk == 32'd2766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	916   :   assert (rdbk == 32'd9797) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	917   :   assert (rdbk == 32'd1021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	918   :   assert (rdbk == 32'd7320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	919   :   assert (rdbk == 32'd3460) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	920   :   assert (rdbk == 32'd5849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	921   :   assert (rdbk == 32'd4764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	922   :   assert (rdbk == 32'd4496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	923   :   assert (rdbk == 32'd1590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	924   :   assert (rdbk == 32'd10785) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	925   :   assert (rdbk == 32'd7963) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	926   :   assert (rdbk == 32'd9156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	927   :   assert (rdbk == 32'd3823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	928   :   assert (rdbk == 32'd8440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	929   :   assert (rdbk == 32'd7431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	930   :   assert (rdbk == 32'd11985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	931   :   assert (rdbk == 32'd1813) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	932   :   assert (rdbk == 32'd8294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	933   :   assert (rdbk == 32'd333) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	934   :   assert (rdbk == 32'd2819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	935   :   assert (rdbk == 32'd1315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	936   :   assert (rdbk == 32'd5125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	937   :   assert (rdbk == 32'd10219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	938   :   assert (rdbk == 32'd3029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	939   :   assert (rdbk == 32'd1021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	940   :   assert (rdbk == 32'd1107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	941   :   assert (rdbk == 32'd4023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	942   :   assert (rdbk == 32'd10019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	943   :   assert (rdbk == 32'd12223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	944   :   assert (rdbk == 32'd6310) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	945   :   assert (rdbk == 32'd12054) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	946   :   assert (rdbk == 32'd7680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	947   :   assert (rdbk == 32'd10999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	948   :   assert (rdbk == 32'd7734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	949   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	950   :   assert (rdbk == 32'd2587) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	951   :   assert (rdbk == 32'd680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	952   :   assert (rdbk == 32'd3000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	953   :   assert (rdbk == 32'd4632) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	954   :   assert (rdbk == 32'd8608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	955   :   assert (rdbk == 32'd8859) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	956   :   assert (rdbk == 32'd2429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	957   :   assert (rdbk == 32'd11232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	958   :   assert (rdbk == 32'd2622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	959   :   assert (rdbk == 32'd6641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	960   :   assert (rdbk == 32'd4520) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	961   :   assert (rdbk == 32'd9522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	962   :   assert (rdbk == 32'd4442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	963   :   assert (rdbk == 32'd7312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	964   :   assert (rdbk == 32'd3089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	965   :   assert (rdbk == 32'd7560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	966   :   assert (rdbk == 32'd10622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	967   :   assert (rdbk == 32'd6280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	968   :   assert (rdbk == 32'd5464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	969   :   assert (rdbk == 32'd4180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	970   :   assert (rdbk == 32'd7974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	971   :   assert (rdbk == 32'd2365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	972   :   assert (rdbk == 32'd2414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	973   :   assert (rdbk == 32'd872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	974   :   assert (rdbk == 32'd656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	975   :   assert (rdbk == 32'd8956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	976   :   assert (rdbk == 32'd6630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	977   :   assert (rdbk == 32'd8287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	978   :   assert (rdbk == 32'd10527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	979   :   assert (rdbk == 32'd11047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	980   :   assert (rdbk == 32'd4752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	981   :   assert (rdbk == 32'd8244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	982   :   assert (rdbk == 32'd9886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	983   :   assert (rdbk == 32'd4409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	984   :   assert (rdbk == 32'd2404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	985   :   assert (rdbk == 32'd12024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	986   :   assert (rdbk == 32'd1892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	987   :   assert (rdbk == 32'd8732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	988   :   assert (rdbk == 32'd2897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	989   :   assert (rdbk == 32'd4841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	990   :   assert (rdbk == 32'd4950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	991   :   assert (rdbk == 32'd12236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	992   :   assert (rdbk == 32'd6976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	993   :   assert (rdbk == 32'd2983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	994   :   assert (rdbk == 32'd2006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	995   :   assert (rdbk == 32'd11065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	996   :   assert (rdbk == 32'd9029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	997   :   assert (rdbk == 32'd4067) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	998   :   assert (rdbk == 32'd3719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	999   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1000   :   assert (rdbk == 32'd5194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1001   :   assert (rdbk == 32'd7619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1002   :   assert (rdbk == 32'd2080) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1003   :   assert (rdbk == 32'd8898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1004   :   assert (rdbk == 32'd2821) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1005   :   assert (rdbk == 32'd6363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1006   :   assert (rdbk == 32'd5697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1007   :   assert (rdbk == 32'd3777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1008   :   assert (rdbk == 32'd9416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1009   :   assert (rdbk == 32'd534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1010   :   assert (rdbk == 32'd9793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1011   :   assert (rdbk == 32'd9051) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1012   :   assert (rdbk == 32'd6480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1013   :   assert (rdbk == 32'd7324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1014   :   assert (rdbk == 32'd11620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1015   :   assert (rdbk == 32'd7411) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1016   :   assert (rdbk == 32'd11198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1017   :   assert (rdbk == 32'd1298) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1018   :   assert (rdbk == 32'd1011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1019   :   assert (rdbk == 32'd10767) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1020   :   assert (rdbk == 32'd10026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1021   :   assert (rdbk == 32'd4756) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1022   :   assert (rdbk == 32'd3028) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1023   :   assert (rdbk == 32'd4733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
    endcase
end

