// Copyright Copyright Fraunhofer Institute for Applied and Integrated Security (AISEC).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

  $fwrite(f,"----------------------------------------------------------------\n");   
  $fwrite(f,"-- PQ-POLY_UNIFORM \n");
  $fwrite(f,"----------------------------------------------------------------\n");   
     
  // Write IMEM from File
  write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq_expand_a.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

  $fwrite(f,"-- IMEM\n");
  // Read IMEM  
  for (int i=0 ; i<129 ; i++) begin 
      //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
  end     

   // Write DMEM from File
  write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq_expand_a.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

  $fwrite(f,"-- DMEM\n");
  // Read DMEM  
  for (int i=0 ; i<16 ; i++) begin 
      //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
  end   
	   
  $fwrite(f,"----------------------------------------------------------------\n");   

  // Set Instruction Counter to zero (optional)
  write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );

  // Start Programm in IMEM
  write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(CmdExecute), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
  cc_start = cc;
  // Poll on Status Register until Programm is finished
  rdbk = '1;
  while (rdbk != '0) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
  end 

  // Measure CC
  cc_stop = cc; 
  cc_count_poly_uniform = cc_stop - cc_start;        
       
  // Read DMEM  
  for (int i=0 ; i<4096 ; i++) begin 
    read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+1024), .tl_o(tl_o), .tl_i(tl_i_d) );
    case(i)
	0   :   assert (rdbk == 32'h163f56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1   :   assert (rdbk == 32'hd88cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2   :   assert (rdbk == 32'h68a78f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3   :   assert (rdbk == 32'h2510fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4   :   assert (rdbk == 32'h30ef1f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	5   :   assert (rdbk == 32'h4e5d23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	6   :   assert (rdbk == 32'h142ef6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	7   :   assert (rdbk == 32'h65db46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	8   :   assert (rdbk == 32'h34304b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	9   :   assert (rdbk == 32'h7877d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	10   :   assert (rdbk == 32'h1bd4c4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	11   :   assert (rdbk == 32'h1ace6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	12   :   assert (rdbk == 32'h46f751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	13   :   assert (rdbk == 32'h607b2a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	14   :   assert (rdbk == 32'h18568e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	15   :   assert (rdbk == 32'h35415f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	16   :   assert (rdbk == 32'h3930da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	17   :   assert (rdbk == 32'h7006e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	18   :   assert (rdbk == 32'h25fa4e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	19   :   assert (rdbk == 32'h556733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	20   :   assert (rdbk == 32'h38a8fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	21   :   assert (rdbk == 32'h2662f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	22   :   assert (rdbk == 32'ha3aad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	23   :   assert (rdbk == 32'h78f859) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	24   :   assert (rdbk == 32'h19b7c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	25   :   assert (rdbk == 32'h46f38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	26   :   assert (rdbk == 32'h7bb802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	27   :   assert (rdbk == 32'h1932b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	28   :   assert (rdbk == 32'h22dd24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	29   :   assert (rdbk == 32'h6eba9e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	30   :   assert (rdbk == 32'h274d3c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	31   :   assert (rdbk == 32'h322d40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	32   :   assert (rdbk == 32'h464435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	33   :   assert (rdbk == 32'h1823e6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	34   :   assert (rdbk == 32'h38e751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	35   :   assert (rdbk == 32'h73bf6a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	36   :   assert (rdbk == 32'h20c953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	37   :   assert (rdbk == 32'h69a5b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	38   :   assert (rdbk == 32'h1d385c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	39   :   assert (rdbk == 32'h32316d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	40   :   assert (rdbk == 32'h157e78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	41   :   assert (rdbk == 32'h6adf19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	42   :   assert (rdbk == 32'h583dee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	43   :   assert (rdbk == 32'h75565e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	44   :   assert (rdbk == 32'h2c6816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	45   :   assert (rdbk == 32'h77d832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	46   :   assert (rdbk == 32'h18db17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	47   :   assert (rdbk == 32'h3304b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	48   :   assert (rdbk == 32'h6bf6f9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	49   :   assert (rdbk == 32'h2ca1a9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	50   :   assert (rdbk == 32'h2725f4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	51   :   assert (rdbk == 32'h1879ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	52   :   assert (rdbk == 32'h4c493e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	53   :   assert (rdbk == 32'h2d890c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	54   :   assert (rdbk == 32'h30bd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	55   :   assert (rdbk == 32'h1579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	56   :   assert (rdbk == 32'h6426e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	57   :   assert (rdbk == 32'h7f80f4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	58   :   assert (rdbk == 32'h3d3a63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	59   :   assert (rdbk == 32'hbaff7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	60   :   assert (rdbk == 32'h624727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	61   :   assert (rdbk == 32'h63ea6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	62   :   assert (rdbk == 32'h3ccc71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	63   :   assert (rdbk == 32'h7c8021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	64   :   assert (rdbk == 32'h3519fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	65   :   assert (rdbk == 32'h5c845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	66   :   assert (rdbk == 32'h509f73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	67   :   assert (rdbk == 32'h5c12fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	68   :   assert (rdbk == 32'h2ab7ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	69   :   assert (rdbk == 32'h58eaac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	70   :   assert (rdbk == 32'h677230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	71   :   assert (rdbk == 32'h3fffc8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	72   :   assert (rdbk == 32'h3e0145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	73   :   assert (rdbk == 32'h5c78b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	74   :   assert (rdbk == 32'h6a0f0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	75   :   assert (rdbk == 32'h1207de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	76   :   assert (rdbk == 32'h5f20db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	77   :   assert (rdbk == 32'h2136c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	78   :   assert (rdbk == 32'h442d89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	79   :   assert (rdbk == 32'h25656c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	80   :   assert (rdbk == 32'h6de7c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	81   :   assert (rdbk == 32'hc499a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	82   :   assert (rdbk == 32'h259422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	83   :   assert (rdbk == 32'h88bd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	84   :   assert (rdbk == 32'hdba25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	85   :   assert (rdbk == 32'h8df83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	86   :   assert (rdbk == 32'hb6e48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	87   :   assert (rdbk == 32'h504653) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	88   :   assert (rdbk == 32'h3e3bbd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	89   :   assert (rdbk == 32'h32f1df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	90   :   assert (rdbk == 32'h6e256b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	91   :   assert (rdbk == 32'h4caeda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	92   :   assert (rdbk == 32'h5cef61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	93   :   assert (rdbk == 32'h331929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	94   :   assert (rdbk == 32'h22eb57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	95   :   assert (rdbk == 32'h5b000d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	96   :   assert (rdbk == 32'h505c6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	97   :   assert (rdbk == 32'h3c6ea4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	98   :   assert (rdbk == 32'h3c0b12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	99   :   assert (rdbk == 32'h272958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	100   :   assert (rdbk == 32'h6fa4d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	101   :   assert (rdbk == 32'h6cf330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	102   :   assert (rdbk == 32'h5ec16e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	103   :   assert (rdbk == 32'h51ad91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	104   :   assert (rdbk == 32'h2d4538) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	105   :   assert (rdbk == 32'he4da9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	106   :   assert (rdbk == 32'h257b43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	107   :   assert (rdbk == 32'h6ad8e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	108   :   assert (rdbk == 32'h2df1fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	109   :   assert (rdbk == 32'h2857) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	110   :   assert (rdbk == 32'h39be2d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	111   :   assert (rdbk == 32'h1d19a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	112   :   assert (rdbk == 32'h25366f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	113   :   assert (rdbk == 32'h11743d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	114   :   assert (rdbk == 32'h6464f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	115   :   assert (rdbk == 32'h7406ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	116   :   assert (rdbk == 32'h934db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	117   :   assert (rdbk == 32'h2480f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	118   :   assert (rdbk == 32'h53f16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	119   :   assert (rdbk == 32'h4b69ef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	120   :   assert (rdbk == 32'h6a5f8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	121   :   assert (rdbk == 32'h703e59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	122   :   assert (rdbk == 32'h575b99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	123   :   assert (rdbk == 32'h1c21d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	124   :   assert (rdbk == 32'h216e4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	125   :   assert (rdbk == 32'h1f8e6d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	126   :   assert (rdbk == 32'h1f537c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	127   :   assert (rdbk == 32'h76975f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	128   :   assert (rdbk == 32'h6bb334) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	129   :   assert (rdbk == 32'h5e6d39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	130   :   assert (rdbk == 32'h5aee28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	131   :   assert (rdbk == 32'h4351ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	132   :   assert (rdbk == 32'h276df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	133   :   assert (rdbk == 32'h72c1cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	134   :   assert (rdbk == 32'h6bd069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	135   :   assert (rdbk == 32'h446546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	136   :   assert (rdbk == 32'h32b5fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	137   :   assert (rdbk == 32'h684a2a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	138   :   assert (rdbk == 32'h75fd8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	139   :   assert (rdbk == 32'h63a74b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	140   :   assert (rdbk == 32'h78adf8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	141   :   assert (rdbk == 32'h5257ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	142   :   assert (rdbk == 32'h19a364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	143   :   assert (rdbk == 32'h728f51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	144   :   assert (rdbk == 32'h631a22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	145   :   assert (rdbk == 32'h62ae01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	146   :   assert (rdbk == 32'h602c17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	147   :   assert (rdbk == 32'h367ca0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	148   :   assert (rdbk == 32'h4abc30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	149   :   assert (rdbk == 32'he1aa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	150   :   assert (rdbk == 32'h5bbe90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	151   :   assert (rdbk == 32'h554357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	152   :   assert (rdbk == 32'h7640a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	153   :   assert (rdbk == 32'h28ae01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	154   :   assert (rdbk == 32'h44c65f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	155   :   assert (rdbk == 32'h6b8ef8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	156   :   assert (rdbk == 32'h6052ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	157   :   assert (rdbk == 32'h6300c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	158   :   assert (rdbk == 32'h374bb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	159   :   assert (rdbk == 32'h282a15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	160   :   assert (rdbk == 32'h440cd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	161   :   assert (rdbk == 32'h68e157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	162   :   assert (rdbk == 32'h1eaae9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	163   :   assert (rdbk == 32'h338c53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	164   :   assert (rdbk == 32'h2e29f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	165   :   assert (rdbk == 32'h2332e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	166   :   assert (rdbk == 32'h7ed1b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	167   :   assert (rdbk == 32'h419826) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	168   :   assert (rdbk == 32'h7b30d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	169   :   assert (rdbk == 32'h68a20a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	170   :   assert (rdbk == 32'h4abd9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	171   :   assert (rdbk == 32'h1c2170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	172   :   assert (rdbk == 32'h12b7af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	173   :   assert (rdbk == 32'h489001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	174   :   assert (rdbk == 32'h35e95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	175   :   assert (rdbk == 32'h624674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	176   :   assert (rdbk == 32'h3290f4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	177   :   assert (rdbk == 32'h7d6af0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	178   :   assert (rdbk == 32'hf1344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	179   :   assert (rdbk == 32'h33ca4f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	180   :   assert (rdbk == 32'h3acd03) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	181   :   assert (rdbk == 32'h17f0e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	182   :   assert (rdbk == 32'h1e7937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	183   :   assert (rdbk == 32'h75e11b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	184   :   assert (rdbk == 32'h7c7936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	185   :   assert (rdbk == 32'h75511e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	186   :   assert (rdbk == 32'h1aa7ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	187   :   assert (rdbk == 32'h258582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	188   :   assert (rdbk == 32'h5a91aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	189   :   assert (rdbk == 32'h1f17f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	190   :   assert (rdbk == 32'h12acb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	191   :   assert (rdbk == 32'h3258bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	192   :   assert (rdbk == 32'h60a93d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	193   :   assert (rdbk == 32'h68905a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	194   :   assert (rdbk == 32'h495d60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	195   :   assert (rdbk == 32'h58c9d9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	196   :   assert (rdbk == 32'h87b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	197   :   assert (rdbk == 32'h591ed1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	198   :   assert (rdbk == 32'h66dcb0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	199   :   assert (rdbk == 32'hb87c4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	200   :   assert (rdbk == 32'hefa5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	201   :   assert (rdbk == 32'hf89ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	202   :   assert (rdbk == 32'h4a352c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	203   :   assert (rdbk == 32'h709d29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	204   :   assert (rdbk == 32'h58b090) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	205   :   assert (rdbk == 32'h5cb571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	206   :   assert (rdbk == 32'h4106f9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	207   :   assert (rdbk == 32'h6963a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	208   :   assert (rdbk == 32'h6c3077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	209   :   assert (rdbk == 32'h4144a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	210   :   assert (rdbk == 32'h4a2997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	211   :   assert (rdbk == 32'h447564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	212   :   assert (rdbk == 32'h3d112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	213   :   assert (rdbk == 32'hc49a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	214   :   assert (rdbk == 32'h52ca2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	215   :   assert (rdbk == 32'h1edddd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	216   :   assert (rdbk == 32'h418d04) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	217   :   assert (rdbk == 32'h2398b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	218   :   assert (rdbk == 32'h3d4b35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	219   :   assert (rdbk == 32'h183f04) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	220   :   assert (rdbk == 32'hbe85f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	221   :   assert (rdbk == 32'h778ba4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	222   :   assert (rdbk == 32'h5255bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	223   :   assert (rdbk == 32'h73fc8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	224   :   assert (rdbk == 32'h49c67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	225   :   assert (rdbk == 32'h14b214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	226   :   assert (rdbk == 32'h5479c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	227   :   assert (rdbk == 32'h5ae529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	228   :   assert (rdbk == 32'h57e08e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	229   :   assert (rdbk == 32'h1ee6bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	230   :   assert (rdbk == 32'h6730ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	231   :   assert (rdbk == 32'h1c5dc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	232   :   assert (rdbk == 32'h759eb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	233   :   assert (rdbk == 32'h67d494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	234   :   assert (rdbk == 32'h19dc0e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	235   :   assert (rdbk == 32'h9a6a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	236   :   assert (rdbk == 32'h2d4f85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	237   :   assert (rdbk == 32'h154b9d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	238   :   assert (rdbk == 32'h507b9d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	239   :   assert (rdbk == 32'h1248b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	240   :   assert (rdbk == 32'h2ca815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	241   :   assert (rdbk == 32'h1a01b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	242   :   assert (rdbk == 32'h464da8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	243   :   assert (rdbk == 32'h35b439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	244   :   assert (rdbk == 32'h6ef866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	245   :   assert (rdbk == 32'h34c54a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	246   :   assert (rdbk == 32'h16b805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	247   :   assert (rdbk == 32'h7d893a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	248   :   assert (rdbk == 32'h2c8fa7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	249   :   assert (rdbk == 32'h52f6c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	250   :   assert (rdbk == 32'h8b150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	251   :   assert (rdbk == 32'h3a40e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	252   :   assert (rdbk == 32'h8923e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	253   :   assert (rdbk == 32'h34f89a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	254   :   assert (rdbk == 32'h1e212c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	255   :   assert (rdbk == 32'h510308) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h1
	256   :   assert (rdbk == 32'hc2f81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	257   :   assert (rdbk == 32'h13710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	258   :   assert (rdbk == 32'h57b6de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	259   :   assert (rdbk == 32'h624a13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	260   :   assert (rdbk == 32'h5e99ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	261   :   assert (rdbk == 32'h4eb5e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	262   :   assert (rdbk == 32'h6880f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	263   :   assert (rdbk == 32'h74997d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	264   :   assert (rdbk == 32'h57a9ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	265   :   assert (rdbk == 32'hf566f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	266   :   assert (rdbk == 32'h45fc01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	267   :   assert (rdbk == 32'h3e2c54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	268   :   assert (rdbk == 32'h7cee0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	269   :   assert (rdbk == 32'h55671) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	270   :   assert (rdbk == 32'h19cce5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	271   :   assert (rdbk == 32'h6d6241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	272   :   assert (rdbk == 32'h10361e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	273   :   assert (rdbk == 32'h61c797) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	274   :   assert (rdbk == 32'h12426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	275   :   assert (rdbk == 32'hfa163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	276   :   assert (rdbk == 32'h181ed4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	277   :   assert (rdbk == 32'h437406) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	278   :   assert (rdbk == 32'h3784ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	279   :   assert (rdbk == 32'h634788) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	280   :   assert (rdbk == 32'h6943ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	281   :   assert (rdbk == 32'h35c2fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	282   :   assert (rdbk == 32'h522d53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	283   :   assert (rdbk == 32'h333914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	284   :   assert (rdbk == 32'h434554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	285   :   assert (rdbk == 32'h35eb98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	286   :   assert (rdbk == 32'h77ae76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	287   :   assert (rdbk == 32'h1363bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	288   :   assert (rdbk == 32'h34de22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	289   :   assert (rdbk == 32'h17046b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	290   :   assert (rdbk == 32'h491c3b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	291   :   assert (rdbk == 32'h58b27a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	292   :   assert (rdbk == 32'h3b38fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	293   :   assert (rdbk == 32'h3c0140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	294   :   assert (rdbk == 32'h3e015d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	295   :   assert (rdbk == 32'h565059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	296   :   assert (rdbk == 32'h207c80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	297   :   assert (rdbk == 32'h4a1e26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	298   :   assert (rdbk == 32'h5f51d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	299   :   assert (rdbk == 32'h1c9ded) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	300   :   assert (rdbk == 32'h2c3b1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	301   :   assert (rdbk == 32'h416e35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	302   :   assert (rdbk == 32'h323622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	303   :   assert (rdbk == 32'h247884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	304   :   assert (rdbk == 32'h6d52ec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	305   :   assert (rdbk == 32'h15b1ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	306   :   assert (rdbk == 32'h15ee74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	307   :   assert (rdbk == 32'h38a322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	308   :   assert (rdbk == 32'h6fecc4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	309   :   assert (rdbk == 32'h33abad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	310   :   assert (rdbk == 32'h32dee2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	311   :   assert (rdbk == 32'h124647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	312   :   assert (rdbk == 32'h271c7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	313   :   assert (rdbk == 32'h1d8b32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	314   :   assert (rdbk == 32'h97aa0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	315   :   assert (rdbk == 32'h1e56c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	316   :   assert (rdbk == 32'h44e157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	317   :   assert (rdbk == 32'h479e00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	318   :   assert (rdbk == 32'h61fffa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	319   :   assert (rdbk == 32'h3fb55f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	320   :   assert (rdbk == 32'h59df1d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	321   :   assert (rdbk == 32'h1a84d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	322   :   assert (rdbk == 32'h73f27b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	323   :   assert (rdbk == 32'h11e3b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	324   :   assert (rdbk == 32'h1f7d91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	325   :   assert (rdbk == 32'h5db8ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	326   :   assert (rdbk == 32'h5110f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	327   :   assert (rdbk == 32'h398307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	328   :   assert (rdbk == 32'h6666e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	329   :   assert (rdbk == 32'h47f9ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	330   :   assert (rdbk == 32'h4f39b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	331   :   assert (rdbk == 32'h22526d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	332   :   assert (rdbk == 32'h4413ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	333   :   assert (rdbk == 32'h1c4d94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	334   :   assert (rdbk == 32'h3bc0ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	335   :   assert (rdbk == 32'h3c8677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	336   :   assert (rdbk == 32'h7234b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	337   :   assert (rdbk == 32'h5d4392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	338   :   assert (rdbk == 32'h710e2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	339   :   assert (rdbk == 32'h67b3f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	340   :   assert (rdbk == 32'h377e34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	341   :   assert (rdbk == 32'h1e2970) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	342   :   assert (rdbk == 32'h24a493) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	343   :   assert (rdbk == 32'h6750d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	344   :   assert (rdbk == 32'h7d5eae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	345   :   assert (rdbk == 32'h72a3d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	346   :   assert (rdbk == 32'h44dcfe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	347   :   assert (rdbk == 32'h2ada35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	348   :   assert (rdbk == 32'h9d7aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	349   :   assert (rdbk == 32'h575c11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	350   :   assert (rdbk == 32'h12eb5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	351   :   assert (rdbk == 32'h7467d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	352   :   assert (rdbk == 32'h43466d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	353   :   assert (rdbk == 32'h37b152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	354   :   assert (rdbk == 32'h7ed208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	355   :   assert (rdbk == 32'h2d0f11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	356   :   assert (rdbk == 32'h4c5fb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	357   :   assert (rdbk == 32'h5a2d65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	358   :   assert (rdbk == 32'h6500ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	359   :   assert (rdbk == 32'h1f6d8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	360   :   assert (rdbk == 32'h22c58f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	361   :   assert (rdbk == 32'h762087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	362   :   assert (rdbk == 32'h98b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	363   :   assert (rdbk == 32'h632a36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	364   :   assert (rdbk == 32'h44548b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	365   :   assert (rdbk == 32'h1c2871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	366   :   assert (rdbk == 32'h38b481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	367   :   assert (rdbk == 32'h21cead) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	368   :   assert (rdbk == 32'ha016b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	369   :   assert (rdbk == 32'h1f18c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	370   :   assert (rdbk == 32'h2118a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	371   :   assert (rdbk == 32'h17710a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	372   :   assert (rdbk == 32'h54a363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	373   :   assert (rdbk == 32'h7694fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	374   :   assert (rdbk == 32'h483ec2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	375   :   assert (rdbk == 32'h160417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	376   :   assert (rdbk == 32'h230aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	377   :   assert (rdbk == 32'h17f673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	378   :   assert (rdbk == 32'h50479c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	379   :   assert (rdbk == 32'h14fd8d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	380   :   assert (rdbk == 32'h135db9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	381   :   assert (rdbk == 32'h6b6d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	382   :   assert (rdbk == 32'h2b8af4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	383   :   assert (rdbk == 32'hd4d6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	384   :   assert (rdbk == 32'h17494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	385   :   assert (rdbk == 32'h63a891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	386   :   assert (rdbk == 32'h475acb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	387   :   assert (rdbk == 32'h53bac7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	388   :   assert (rdbk == 32'h365723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	389   :   assert (rdbk == 32'h18f6c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	390   :   assert (rdbk == 32'h4c7acb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	391   :   assert (rdbk == 32'h200e0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	392   :   assert (rdbk == 32'h5f15cd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	393   :   assert (rdbk == 32'h42cbef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	394   :   assert (rdbk == 32'h77351e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	395   :   assert (rdbk == 32'h59777f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	396   :   assert (rdbk == 32'h114693) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	397   :   assert (rdbk == 32'h78d492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	398   :   assert (rdbk == 32'h6810bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	399   :   assert (rdbk == 32'h3b14af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	400   :   assert (rdbk == 32'h3a344c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	401   :   assert (rdbk == 32'h5e592f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	402   :   assert (rdbk == 32'h262a1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	403   :   assert (rdbk == 32'h50d656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	404   :   assert (rdbk == 32'h30ce0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	405   :   assert (rdbk == 32'h140441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	406   :   assert (rdbk == 32'h180790) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	407   :   assert (rdbk == 32'h777c3e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	408   :   assert (rdbk == 32'h288d71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	409   :   assert (rdbk == 32'h3e1de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	410   :   assert (rdbk == 32'h69a0f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	411   :   assert (rdbk == 32'h52d18d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	412   :   assert (rdbk == 32'h1a1a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	413   :   assert (rdbk == 32'h6e6774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	414   :   assert (rdbk == 32'h336a04) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	415   :   assert (rdbk == 32'h196a19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	416   :   assert (rdbk == 32'h1c0004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	417   :   assert (rdbk == 32'h11c60d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	418   :   assert (rdbk == 32'h4a3392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	419   :   assert (rdbk == 32'h334be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	420   :   assert (rdbk == 32'h4f3f82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	421   :   assert (rdbk == 32'h1339d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	422   :   assert (rdbk == 32'h148040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	423   :   assert (rdbk == 32'h133bcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	424   :   assert (rdbk == 32'h47ed4d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	425   :   assert (rdbk == 32'h11b5a1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	426   :   assert (rdbk == 32'h175525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	427   :   assert (rdbk == 32'h2c18ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	428   :   assert (rdbk == 32'h7bfe4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	429   :   assert (rdbk == 32'h499d8e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	430   :   assert (rdbk == 32'h449b50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	431   :   assert (rdbk == 32'h7d4d53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	432   :   assert (rdbk == 32'h5ac240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	433   :   assert (rdbk == 32'h350736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	434   :   assert (rdbk == 32'h66a432) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	435   :   assert (rdbk == 32'h6f9d38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	436   :   assert (rdbk == 32'h6131fe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	437   :   assert (rdbk == 32'h97b55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	438   :   assert (rdbk == 32'h5f207b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	439   :   assert (rdbk == 32'h20cc2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	440   :   assert (rdbk == 32'h11088e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	441   :   assert (rdbk == 32'h315581) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	442   :   assert (rdbk == 32'h30416e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	443   :   assert (rdbk == 32'h416f3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	444   :   assert (rdbk == 32'h7b65a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	445   :   assert (rdbk == 32'h34aa3e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	446   :   assert (rdbk == 32'he99cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	447   :   assert (rdbk == 32'h6b26ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	448   :   assert (rdbk == 32'hfee87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	449   :   assert (rdbk == 32'h20aabd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	450   :   assert (rdbk == 32'h58a2eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	451   :   assert (rdbk == 32'h40c67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	452   :   assert (rdbk == 32'h3945b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	453   :   assert (rdbk == 32'h7f7325) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	454   :   assert (rdbk == 32'h527b83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	455   :   assert (rdbk == 32'h148765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	456   :   assert (rdbk == 32'h2e8f0c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	457   :   assert (rdbk == 32'h56a780) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	458   :   assert (rdbk == 32'h6496e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	459   :   assert (rdbk == 32'h71a71a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	460   :   assert (rdbk == 32'h53bf8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	461   :   assert (rdbk == 32'h39cf41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	462   :   assert (rdbk == 32'h7294ae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	463   :   assert (rdbk == 32'h5d3881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	464   :   assert (rdbk == 32'h43f761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	465   :   assert (rdbk == 32'he8699) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	466   :   assert (rdbk == 32'h271b5e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	467   :   assert (rdbk == 32'h65383f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	468   :   assert (rdbk == 32'h52fee5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	469   :   assert (rdbk == 32'h20ed23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	470   :   assert (rdbk == 32'h4770fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	471   :   assert (rdbk == 32'h166f43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	472   :   assert (rdbk == 32'h64741c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	473   :   assert (rdbk == 32'h2ad914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	474   :   assert (rdbk == 32'h23a09e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	475   :   assert (rdbk == 32'h105097) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	476   :   assert (rdbk == 32'h119fb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	477   :   assert (rdbk == 32'h18ad63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	478   :   assert (rdbk == 32'h44fa00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	479   :   assert (rdbk == 32'h31815c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	480   :   assert (rdbk == 32'hc0a57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	481   :   assert (rdbk == 32'h8fdaf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	482   :   assert (rdbk == 32'h3a70fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	483   :   assert (rdbk == 32'h712e74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	484   :   assert (rdbk == 32'h4d5ec0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	485   :   assert (rdbk == 32'h35ed9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	486   :   assert (rdbk == 32'h114a83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	487   :   assert (rdbk == 32'hf81da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	488   :   assert (rdbk == 32'h1f7d7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	489   :   assert (rdbk == 32'h4d3db1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	490   :   assert (rdbk == 32'h1367de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	491   :   assert (rdbk == 32'h62fb5c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	492   :   assert (rdbk == 32'h2d0279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	493   :   assert (rdbk == 32'h7987ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	494   :   assert (rdbk == 32'h25a3b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	495   :   assert (rdbk == 32'h486234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	496   :   assert (rdbk == 32'h229b2a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	497   :   assert (rdbk == 32'h43a0e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	498   :   assert (rdbk == 32'hd13af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	499   :   assert (rdbk == 32'h786494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	500   :   assert (rdbk == 32'h5fcf77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	501   :   assert (rdbk == 32'h63673f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	502   :   assert (rdbk == 32'h59a343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	503   :   assert (rdbk == 32'h4d1d9e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	504   :   assert (rdbk == 32'h5fae60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	505   :   assert (rdbk == 32'h100f64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	506   :   assert (rdbk == 32'h236f55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	507   :   assert (rdbk == 32'h2e68c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	508   :   assert (rdbk == 32'h4ad2ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	509   :   assert (rdbk == 32'h16bb93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	510   :   assert (rdbk == 32'h5e071c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	511   :   assert (rdbk == 32'h76f79e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h2
	512   :   assert (rdbk == 32'h22aea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	513   :   assert (rdbk == 32'h7453bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	514   :   assert (rdbk == 32'h581f87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	515   :   assert (rdbk == 32'h7b54b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	516   :   assert (rdbk == 32'h321e7c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	517   :   assert (rdbk == 32'h24ecf9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	518   :   assert (rdbk == 32'h2150ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	519   :   assert (rdbk == 32'h697258) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	520   :   assert (rdbk == 32'hd07e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	521   :   assert (rdbk == 32'h1929ec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	522   :   assert (rdbk == 32'h70b877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	523   :   assert (rdbk == 32'h528bcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	524   :   assert (rdbk == 32'hb3d6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	525   :   assert (rdbk == 32'h71331b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	526   :   assert (rdbk == 32'h7f3b5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	527   :   assert (rdbk == 32'h652efe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	528   :   assert (rdbk == 32'h1992bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	529   :   assert (rdbk == 32'h776a96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	530   :   assert (rdbk == 32'h236af3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	531   :   assert (rdbk == 32'h74659d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	532   :   assert (rdbk == 32'h2840f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	533   :   assert (rdbk == 32'h187df9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	534   :   assert (rdbk == 32'he1675) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	535   :   assert (rdbk == 32'h62adf5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	536   :   assert (rdbk == 32'h17ab01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	537   :   assert (rdbk == 32'h610c35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	538   :   assert (rdbk == 32'h2862c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	539   :   assert (rdbk == 32'h5bce45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	540   :   assert (rdbk == 32'h773331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	541   :   assert (rdbk == 32'h137b12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	542   :   assert (rdbk == 32'h55ddb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	543   :   assert (rdbk == 32'h6b5af4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	544   :   assert (rdbk == 32'h306e20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	545   :   assert (rdbk == 32'h12ccd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	546   :   assert (rdbk == 32'h93a0e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	547   :   assert (rdbk == 32'h5c0c84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	548   :   assert (rdbk == 32'h2358c4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	549   :   assert (rdbk == 32'h65ebb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	550   :   assert (rdbk == 32'h3f772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	551   :   assert (rdbk == 32'h2a2769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	552   :   assert (rdbk == 32'h713f60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	553   :   assert (rdbk == 32'h5d611d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	554   :   assert (rdbk == 32'h6c27fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	555   :   assert (rdbk == 32'h28746f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	556   :   assert (rdbk == 32'h365acd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	557   :   assert (rdbk == 32'h77866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	558   :   assert (rdbk == 32'h3de01d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	559   :   assert (rdbk == 32'h16a204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	560   :   assert (rdbk == 32'h1a1df4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	561   :   assert (rdbk == 32'h5c641e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	562   :   assert (rdbk == 32'h10eb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	563   :   assert (rdbk == 32'hf1d03) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	564   :   assert (rdbk == 32'h546207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	565   :   assert (rdbk == 32'h394a2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	566   :   assert (rdbk == 32'h4db37a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	567   :   assert (rdbk == 32'h4803eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	568   :   assert (rdbk == 32'h3da806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	569   :   assert (rdbk == 32'h2a0bca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	570   :   assert (rdbk == 32'h51328f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	571   :   assert (rdbk == 32'h717838) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	572   :   assert (rdbk == 32'h3ced57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	573   :   assert (rdbk == 32'h764d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	574   :   assert (rdbk == 32'h7af6a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	575   :   assert (rdbk == 32'h1e9086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	576   :   assert (rdbk == 32'h455f84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	577   :   assert (rdbk == 32'h1341a9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	578   :   assert (rdbk == 32'h1970ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	579   :   assert (rdbk == 32'h20d850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	580   :   assert (rdbk == 32'h3d26a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	581   :   assert (rdbk == 32'h57a29a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	582   :   assert (rdbk == 32'h4e9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	583   :   assert (rdbk == 32'h5ffcb7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	584   :   assert (rdbk == 32'h6c60bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	585   :   assert (rdbk == 32'h22a2a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	586   :   assert (rdbk == 32'h1c052e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	587   :   assert (rdbk == 32'h355541) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	588   :   assert (rdbk == 32'h1f97b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	589   :   assert (rdbk == 32'h5799c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	590   :   assert (rdbk == 32'h7e4b39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	591   :   assert (rdbk == 32'h333f56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	592   :   assert (rdbk == 32'h15b89d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	593   :   assert (rdbk == 32'h16bbb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	594   :   assert (rdbk == 32'h42322c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	595   :   assert (rdbk == 32'h76bc03) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	596   :   assert (rdbk == 32'h39c477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	597   :   assert (rdbk == 32'h6d616f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	598   :   assert (rdbk == 32'h17b601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	599   :   assert (rdbk == 32'hb3cba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	600   :   assert (rdbk == 32'h425413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	601   :   assert (rdbk == 32'h6908a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	602   :   assert (rdbk == 32'h74abab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	603   :   assert (rdbk == 32'h163484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	604   :   assert (rdbk == 32'h781239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	605   :   assert (rdbk == 32'h173c3d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	606   :   assert (rdbk == 32'h633eb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	607   :   assert (rdbk == 32'h42de39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	608   :   assert (rdbk == 32'h7795b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	609   :   assert (rdbk == 32'h43b601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	610   :   assert (rdbk == 32'h6b434a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	611   :   assert (rdbk == 32'h7c8f98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	612   :   assert (rdbk == 32'h594af4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	613   :   assert (rdbk == 32'h58884c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	614   :   assert (rdbk == 32'h1b92b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	615   :   assert (rdbk == 32'hb4b7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	616   :   assert (rdbk == 32'h7dea7a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	617   :   assert (rdbk == 32'h72ed85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	618   :   assert (rdbk == 32'h751ffb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	619   :   assert (rdbk == 32'h63c29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	620   :   assert (rdbk == 32'h12643d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	621   :   assert (rdbk == 32'h27233a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	622   :   assert (rdbk == 32'h1a850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	623   :   assert (rdbk == 32'h62d120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	624   :   assert (rdbk == 32'h4688f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	625   :   assert (rdbk == 32'h2034f4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	626   :   assert (rdbk == 32'h829b1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	627   :   assert (rdbk == 32'h2ada49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	628   :   assert (rdbk == 32'h786f98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	629   :   assert (rdbk == 32'h561aed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	630   :   assert (rdbk == 32'h2bd30e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	631   :   assert (rdbk == 32'h1a25a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	632   :   assert (rdbk == 32'h4bc7a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	633   :   assert (rdbk == 32'h3cc45e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	634   :   assert (rdbk == 32'h63942d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	635   :   assert (rdbk == 32'h11bf8e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	636   :   assert (rdbk == 32'h4960bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	637   :   assert (rdbk == 32'h591a22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	638   :   assert (rdbk == 32'h438c48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	639   :   assert (rdbk == 32'h179e1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	640   :   assert (rdbk == 32'h566278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	641   :   assert (rdbk == 32'h7a7f89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	642   :   assert (rdbk == 32'h41cbb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	643   :   assert (rdbk == 32'h7031d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	644   :   assert (rdbk == 32'h21e28a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	645   :   assert (rdbk == 32'h5b404e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	646   :   assert (rdbk == 32'h718612) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	647   :   assert (rdbk == 32'h615b67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	648   :   assert (rdbk == 32'h64c342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	649   :   assert (rdbk == 32'h521a12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	650   :   assert (rdbk == 32'h750f18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	651   :   assert (rdbk == 32'h154672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	652   :   assert (rdbk == 32'h11d575) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	653   :   assert (rdbk == 32'h335caf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	654   :   assert (rdbk == 32'h13e9af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	655   :   assert (rdbk == 32'h571188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	656   :   assert (rdbk == 32'h5992aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	657   :   assert (rdbk == 32'h2f903b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	658   :   assert (rdbk == 32'h73adbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	659   :   assert (rdbk == 32'h382d96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	660   :   assert (rdbk == 32'h2f3110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	661   :   assert (rdbk == 32'h1cece2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	662   :   assert (rdbk == 32'h598d4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	663   :   assert (rdbk == 32'h610651) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	664   :   assert (rdbk == 32'h46e61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	665   :   assert (rdbk == 32'h531d18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	666   :   assert (rdbk == 32'h1b49d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	667   :   assert (rdbk == 32'h40168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	668   :   assert (rdbk == 32'h702451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	669   :   assert (rdbk == 32'h2ba5c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	670   :   assert (rdbk == 32'h3bbf36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	671   :   assert (rdbk == 32'h2a40c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	672   :   assert (rdbk == 32'h5d7309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	673   :   assert (rdbk == 32'h5ad30e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	674   :   assert (rdbk == 32'h6a6ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	675   :   assert (rdbk == 32'hc297f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	676   :   assert (rdbk == 32'h23783e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	677   :   assert (rdbk == 32'h92f3f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	678   :   assert (rdbk == 32'h458071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	679   :   assert (rdbk == 32'h1e467a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	680   :   assert (rdbk == 32'h273f90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	681   :   assert (rdbk == 32'h3dfab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	682   :   assert (rdbk == 32'h2f71f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	683   :   assert (rdbk == 32'h6abaa3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	684   :   assert (rdbk == 32'h6c7137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	685   :   assert (rdbk == 32'h576901) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	686   :   assert (rdbk == 32'h22147b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	687   :   assert (rdbk == 32'h22c477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	688   :   assert (rdbk == 32'h4c8a7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	689   :   assert (rdbk == 32'h78937f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	690   :   assert (rdbk == 32'h47567b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	691   :   assert (rdbk == 32'hb6e9c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	692   :   assert (rdbk == 32'h7e7c47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	693   :   assert (rdbk == 32'h780253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	694   :   assert (rdbk == 32'h212bae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	695   :   assert (rdbk == 32'h69c0ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	696   :   assert (rdbk == 32'h17ab4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	697   :   assert (rdbk == 32'h7efcdb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	698   :   assert (rdbk == 32'h63f875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	699   :   assert (rdbk == 32'h1d344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	700   :   assert (rdbk == 32'h369248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	701   :   assert (rdbk == 32'h280e8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	702   :   assert (rdbk == 32'h653dc8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	703   :   assert (rdbk == 32'h227175) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	704   :   assert (rdbk == 32'h53c163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	705   :   assert (rdbk == 32'h10a498) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	706   :   assert (rdbk == 32'h7118f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	707   :   assert (rdbk == 32'h721044) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	708   :   assert (rdbk == 32'h11ea6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	709   :   assert (rdbk == 32'h34750c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	710   :   assert (rdbk == 32'h4cb99f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	711   :   assert (rdbk == 32'h16051e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	712   :   assert (rdbk == 32'h55201b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	713   :   assert (rdbk == 32'hce031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	714   :   assert (rdbk == 32'h43a224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	715   :   assert (rdbk == 32'h7f96ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	716   :   assert (rdbk == 32'h2e5fc5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	717   :   assert (rdbk == 32'h778f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	718   :   assert (rdbk == 32'h37cc15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	719   :   assert (rdbk == 32'h50060c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	720   :   assert (rdbk == 32'h2c3604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	721   :   assert (rdbk == 32'h1b6988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	722   :   assert (rdbk == 32'h58c4cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	723   :   assert (rdbk == 32'h2c8d5c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	724   :   assert (rdbk == 32'h6f5b4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	725   :   assert (rdbk == 32'h4b46cd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	726   :   assert (rdbk == 32'h2d7bbc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	727   :   assert (rdbk == 32'h38f4a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	728   :   assert (rdbk == 32'h37853a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	729   :   assert (rdbk == 32'h4acd54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	730   :   assert (rdbk == 32'h16dbc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	731   :   assert (rdbk == 32'h5ce0b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	732   :   assert (rdbk == 32'h7a4ba2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	733   :   assert (rdbk == 32'h36bc4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	734   :   assert (rdbk == 32'h316c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	735   :   assert (rdbk == 32'h1bbf3c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	736   :   assert (rdbk == 32'h5512c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	737   :   assert (rdbk == 32'h656a12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	738   :   assert (rdbk == 32'h57e969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	739   :   assert (rdbk == 32'h3c0846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	740   :   assert (rdbk == 32'h41cf3c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	741   :   assert (rdbk == 32'hc5117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	742   :   assert (rdbk == 32'h60fb26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	743   :   assert (rdbk == 32'h41e1d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	744   :   assert (rdbk == 32'h4fcb67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	745   :   assert (rdbk == 32'h3dcef3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	746   :   assert (rdbk == 32'h664569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	747   :   assert (rdbk == 32'h376959) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	748   :   assert (rdbk == 32'hd6a4e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	749   :   assert (rdbk == 32'h4352a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	750   :   assert (rdbk == 32'h2549b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	751   :   assert (rdbk == 32'h47b288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	752   :   assert (rdbk == 32'h6e3984) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	753   :   assert (rdbk == 32'h2bf48f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	754   :   assert (rdbk == 32'h14fc99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	755   :   assert (rdbk == 32'h541e0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	756   :   assert (rdbk == 32'h325ca5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	757   :   assert (rdbk == 32'h6d178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	758   :   assert (rdbk == 32'h177841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	759   :   assert (rdbk == 32'h6c8f3f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	760   :   assert (rdbk == 32'h3f669b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	761   :   assert (rdbk == 32'h69e831) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	762   :   assert (rdbk == 32'h31219e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	763   :   assert (rdbk == 32'h26143a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	764   :   assert (rdbk == 32'h4ef54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	765   :   assert (rdbk == 32'h28fc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	766   :   assert (rdbk == 32'h77d3f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	767   :   assert (rdbk == 32'h2b5805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	//Nonce: 32'h3
	768   :   assert (rdbk == 32'h75c2b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	769   :   assert (rdbk == 32'h6ecded) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	770   :   assert (rdbk == 32'h3ad04b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	771   :   assert (rdbk == 32'h18422d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	772   :   assert (rdbk == 32'had66b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	773   :   assert (rdbk == 32'h48674e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	774   :   assert (rdbk == 32'h17e1df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	775   :   assert (rdbk == 32'h7f3864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	776   :   assert (rdbk == 32'h40b2e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	777   :   assert (rdbk == 32'h4c485c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	778   :   assert (rdbk == 32'h364a9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	779   :   assert (rdbk == 32'h3f2a75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	780   :   assert (rdbk == 32'h370016) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	781   :   assert (rdbk == 32'h430ea2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	782   :   assert (rdbk == 32'h21095c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	783   :   assert (rdbk == 32'h45d577) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	784   :   assert (rdbk == 32'h5b97a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	785   :   assert (rdbk == 32'h7d7b56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	786   :   assert (rdbk == 32'h9cb8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	787   :   assert (rdbk == 32'h40fff0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	788   :   assert (rdbk == 32'h6e2cb4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	789   :   assert (rdbk == 32'h71f280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	790   :   assert (rdbk == 32'hc2fef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	791   :   assert (rdbk == 32'h5483cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	792   :   assert (rdbk == 32'h3d4f5e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	793   :   assert (rdbk == 32'h122797) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	794   :   assert (rdbk == 32'h7ad050) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	795   :   assert (rdbk == 32'h32e1a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	796   :   assert (rdbk == 32'h720d95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	797   :   assert (rdbk == 32'h136153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	798   :   assert (rdbk == 32'h378aa1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	799   :   assert (rdbk == 32'h15cf1a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	800   :   assert (rdbk == 32'hb1f4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	801   :   assert (rdbk == 32'h11dd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	802   :   assert (rdbk == 32'h70064e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	803   :   assert (rdbk == 32'h1244d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	804   :   assert (rdbk == 32'hb6042) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	805   :   assert (rdbk == 32'h5a5c76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	806   :   assert (rdbk == 32'h4db02d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	807   :   assert (rdbk == 32'h59c765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	808   :   assert (rdbk == 32'h5399b2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	809   :   assert (rdbk == 32'h6f6513) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	810   :   assert (rdbk == 32'h291373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	811   :   assert (rdbk == 32'h78c50e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	812   :   assert (rdbk == 32'h6140cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	813   :   assert (rdbk == 32'h18e18a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	814   :   assert (rdbk == 32'h401e38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	815   :   assert (rdbk == 32'h7a3cdd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	816   :   assert (rdbk == 32'h18b03) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	817   :   assert (rdbk == 32'h41390c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	818   :   assert (rdbk == 32'h54c1cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	819   :   assert (rdbk == 32'h9e2ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	820   :   assert (rdbk == 32'h12df91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	821   :   assert (rdbk == 32'h17bbf3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	822   :   assert (rdbk == 32'h5527f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	823   :   assert (rdbk == 32'h447b59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	824   :   assert (rdbk == 32'h6379c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	825   :   assert (rdbk == 32'h5c6013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	826   :   assert (rdbk == 32'h2bd80e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	827   :   assert (rdbk == 32'h5c458e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	828   :   assert (rdbk == 32'h3fa060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	829   :   assert (rdbk == 32'h7d3881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	830   :   assert (rdbk == 32'h3b851f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	831   :   assert (rdbk == 32'h6ca883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	832   :   assert (rdbk == 32'h1021f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	833   :   assert (rdbk == 32'h766e1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	834   :   assert (rdbk == 32'h3e7c60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	835   :   assert (rdbk == 32'h6578a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	836   :   assert (rdbk == 32'hd00ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	837   :   assert (rdbk == 32'h11221a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	838   :   assert (rdbk == 32'h7b4397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	839   :   assert (rdbk == 32'h15fb02) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	840   :   assert (rdbk == 32'h21cb0a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	841   :   assert (rdbk == 32'h7d5c7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	842   :   assert (rdbk == 32'h40f4fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	843   :   assert (rdbk == 32'h4db5b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	844   :   assert (rdbk == 32'h4ac3ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	845   :   assert (rdbk == 32'h72308a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	846   :   assert (rdbk == 32'h29af74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	847   :   assert (rdbk == 32'h7e8266) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	848   :   assert (rdbk == 32'h628962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	849   :   assert (rdbk == 32'h5c5c8e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	850   :   assert (rdbk == 32'h11fe6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	851   :   assert (rdbk == 32'h6cf68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	852   :   assert (rdbk == 32'h160654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	853   :   assert (rdbk == 32'h58fed7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	854   :   assert (rdbk == 32'h32aecb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	855   :   assert (rdbk == 32'h5ddd5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	856   :   assert (rdbk == 32'h25824) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	857   :   assert (rdbk == 32'h5d7915) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	858   :   assert (rdbk == 32'hc1a65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	859   :   assert (rdbk == 32'h3e1cc6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	860   :   assert (rdbk == 32'h1f53ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	861   :   assert (rdbk == 32'h222895) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	862   :   assert (rdbk == 32'h626e7b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	863   :   assert (rdbk == 32'h49e3c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	864   :   assert (rdbk == 32'h50936c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	865   :   assert (rdbk == 32'h412f22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	866   :   assert (rdbk == 32'h36abaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	867   :   assert (rdbk == 32'h875e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	868   :   assert (rdbk == 32'h689c6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	869   :   assert (rdbk == 32'h6886c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	870   :   assert (rdbk == 32'h70a30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	871   :   assert (rdbk == 32'h3cbc0a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	872   :   assert (rdbk == 32'h2b9f96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	873   :   assert (rdbk == 32'h694f2e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	874   :   assert (rdbk == 32'h229668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	875   :   assert (rdbk == 32'h546486) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	876   :   assert (rdbk == 32'h5571f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	877   :   assert (rdbk == 32'h5da14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	878   :   assert (rdbk == 32'h69d83b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	879   :   assert (rdbk == 32'h388489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	880   :   assert (rdbk == 32'h3e234a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	881   :   assert (rdbk == 32'h655256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	882   :   assert (rdbk == 32'h276948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	883   :   assert (rdbk == 32'hcaee1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	884   :   assert (rdbk == 32'h274f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	885   :   assert (rdbk == 32'h2e4441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	886   :   assert (rdbk == 32'h1fe766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	887   :   assert (rdbk == 32'h3ba672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	888   :   assert (rdbk == 32'h4c71b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	889   :   assert (rdbk == 32'h5c151a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	890   :   assert (rdbk == 32'h5bc6f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	891   :   assert (rdbk == 32'h384946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	892   :   assert (rdbk == 32'h72f1ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	893   :   assert (rdbk == 32'h6cbb06) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	894   :   assert (rdbk == 32'h548ed3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	895   :   assert (rdbk == 32'h68624c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	896   :   assert (rdbk == 32'h23f047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	897   :   assert (rdbk == 32'h7c018d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	898   :   assert (rdbk == 32'h1309d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	899   :   assert (rdbk == 32'h1abd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	900   :   assert (rdbk == 32'h56c4c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	901   :   assert (rdbk == 32'h1818cd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	902   :   assert (rdbk == 32'h5e66d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	903   :   assert (rdbk == 32'h4c5f06) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	904   :   assert (rdbk == 32'h591041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	905   :   assert (rdbk == 32'h492636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	906   :   assert (rdbk == 32'h21e49f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	907   :   assert (rdbk == 32'h39bbce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	908   :   assert (rdbk == 32'h7241f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	909   :   assert (rdbk == 32'h32e047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	910   :   assert (rdbk == 32'h8319e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	911   :   assert (rdbk == 32'h68e5bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	912   :   assert (rdbk == 32'h4ccef4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	913   :   assert (rdbk == 32'h2e54c6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	914   :   assert (rdbk == 32'h2ff315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	915   :   assert (rdbk == 32'h48ff1e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	916   :   assert (rdbk == 32'h5e86d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	917   :   assert (rdbk == 32'h259285) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	918   :   assert (rdbk == 32'h26c3c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	919   :   assert (rdbk == 32'h344162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	920   :   assert (rdbk == 32'h109f38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	921   :   assert (rdbk == 32'h6329b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	922   :   assert (rdbk == 32'h1ae465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	923   :   assert (rdbk == 32'h518daa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	924   :   assert (rdbk == 32'h6a6b16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	925   :   assert (rdbk == 32'h70b9e1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	926   :   assert (rdbk == 32'h1887fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	927   :   assert (rdbk == 32'h70d8da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	928   :   assert (rdbk == 32'h493ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	929   :   assert (rdbk == 32'h7c719f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	930   :   assert (rdbk == 32'h76d9d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	931   :   assert (rdbk == 32'h47a41c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	932   :   assert (rdbk == 32'h5edf45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	933   :   assert (rdbk == 32'h7eb927) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	934   :   assert (rdbk == 32'h2be0da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	935   :   assert (rdbk == 32'h6af184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	936   :   assert (rdbk == 32'h4eed6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	937   :   assert (rdbk == 32'h412712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	938   :   assert (rdbk == 32'h7fd450) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	939   :   assert (rdbk == 32'h8fcb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	940   :   assert (rdbk == 32'h2e1de0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	941   :   assert (rdbk == 32'h683751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	942   :   assert (rdbk == 32'hea9da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	943   :   assert (rdbk == 32'h3b2c6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	944   :   assert (rdbk == 32'h2a4967) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	945   :   assert (rdbk == 32'h4bc97d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	946   :   assert (rdbk == 32'h13c544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	947   :   assert (rdbk == 32'h7a6c65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	948   :   assert (rdbk == 32'h40d97d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	949   :   assert (rdbk == 32'h71db3c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	950   :   assert (rdbk == 32'h7f51b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	951   :   assert (rdbk == 32'h776c90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	952   :   assert (rdbk == 32'h3f6d02) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	953   :   assert (rdbk == 32'h150f86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	954   :   assert (rdbk == 32'h4830ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	955   :   assert (rdbk == 32'h3ca749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	956   :   assert (rdbk == 32'h259659) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	957   :   assert (rdbk == 32'h5965bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	958   :   assert (rdbk == 32'h261d5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	959   :   assert (rdbk == 32'h489c82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	960   :   assert (rdbk == 32'h6c986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	961   :   assert (rdbk == 32'h6e2b0c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	962   :   assert (rdbk == 32'h37957) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	963   :   assert (rdbk == 32'h60d5a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	964   :   assert (rdbk == 32'h3b60d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	965   :   assert (rdbk == 32'h2e26d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	966   :   assert (rdbk == 32'h25ab89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	967   :   assert (rdbk == 32'h3d3fbe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	968   :   assert (rdbk == 32'h6991b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	969   :   assert (rdbk == 32'h54875b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	970   :   assert (rdbk == 32'h3c45d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	971   :   assert (rdbk == 32'h207d92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	972   :   assert (rdbk == 32'h7b05fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	973   :   assert (rdbk == 32'h3f410b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	974   :   assert (rdbk == 32'h203943) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	975   :   assert (rdbk == 32'h576ab2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	976   :   assert (rdbk == 32'h1adf77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	977   :   assert (rdbk == 32'h6fcb00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	978   :   assert (rdbk == 32'h501ab9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	979   :   assert (rdbk == 32'he6c91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	980   :   assert (rdbk == 32'h483df5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	981   :   assert (rdbk == 32'h698a37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	982   :   assert (rdbk == 32'h7ce856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	983   :   assert (rdbk == 32'h721c27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	984   :   assert (rdbk == 32'h644739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	985   :   assert (rdbk == 32'h5d8fc7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	986   :   assert (rdbk == 32'h44bbbc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	987   :   assert (rdbk == 32'h4c06c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	988   :   assert (rdbk == 32'h2380f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	989   :   assert (rdbk == 32'h752372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	990   :   assert (rdbk == 32'h7c4330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	991   :   assert (rdbk == 32'ha8429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	992   :   assert (rdbk == 32'h69a42a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	993   :   assert (rdbk == 32'h1a9a80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	994   :   assert (rdbk == 32'h1de82f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	995   :   assert (rdbk == 32'h42db71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	996   :   assert (rdbk == 32'h7302eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	997   :   assert (rdbk == 32'h2acabb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	998   :   assert (rdbk == 32'h7e60e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	999   :   assert (rdbk == 32'h6206f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1000   :   assert (rdbk == 32'h44c0e1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1001   :   assert (rdbk == 32'h762a69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1002   :   assert (rdbk == 32'h4a909a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1003   :   assert (rdbk == 32'h17e733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1004   :   assert (rdbk == 32'h616977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1005   :   assert (rdbk == 32'h77c083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1006   :   assert (rdbk == 32'h7f17ae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1007   :   assert (rdbk == 32'h16d418) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1008   :   assert (rdbk == 32'h692c98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1009   :   assert (rdbk == 32'h31fb3b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1010   :   assert (rdbk == 32'h6dda3f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1011   :   assert (rdbk == 32'h780e69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1012   :   assert (rdbk == 32'h413a64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1013   :   assert (rdbk == 32'h6797dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1014   :   assert (rdbk == 32'h3fd8a1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1015   :   assert (rdbk == 32'h3ca355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1016   :   assert (rdbk == 32'h2a3c0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1017   :   assert (rdbk == 32'h54666f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1018   :   assert (rdbk == 32'h73c183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1019   :   assert (rdbk == 32'h3ba78b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1020   :   assert (rdbk == 32'h249264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1021   :   assert (rdbk == 32'h3bfd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1022   :   assert (rdbk == 32'h496197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1023   :   assert (rdbk == 32'h1199f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h100
	1024   :   assert (rdbk == 32'h2cc039) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1025   :   assert (rdbk == 32'h4baff0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1026   :   assert (rdbk == 32'h6cad52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1027   :   assert (rdbk == 32'h83cb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1028   :   assert (rdbk == 32'hadad1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1029   :   assert (rdbk == 32'h48e6fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1030   :   assert (rdbk == 32'h364b53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1031   :   assert (rdbk == 32'h116fda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1032   :   assert (rdbk == 32'h2becf8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1033   :   assert (rdbk == 32'h401b65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1034   :   assert (rdbk == 32'hdc456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1035   :   assert (rdbk == 32'h3ebebe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1036   :   assert (rdbk == 32'h791c88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1037   :   assert (rdbk == 32'h266e59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1038   :   assert (rdbk == 32'h5e37ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1039   :   assert (rdbk == 32'h5ee4b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1040   :   assert (rdbk == 32'h230863) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1041   :   assert (rdbk == 32'h71e45c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1042   :   assert (rdbk == 32'h7220da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1043   :   assert (rdbk == 32'h486bc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1044   :   assert (rdbk == 32'h31dc9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1045   :   assert (rdbk == 32'h542b03) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1046   :   assert (rdbk == 32'h77b020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1047   :   assert (rdbk == 32'h6effdd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1048   :   assert (rdbk == 32'h60e6b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1049   :   assert (rdbk == 32'h72bd5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1050   :   assert (rdbk == 32'h1de8f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1051   :   assert (rdbk == 32'hc7947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1052   :   assert (rdbk == 32'h5f910d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1053   :   assert (rdbk == 32'h3a8a17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1054   :   assert (rdbk == 32'h7b3e63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1055   :   assert (rdbk == 32'h142564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1056   :   assert (rdbk == 32'h1050b1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1057   :   assert (rdbk == 32'h20edf5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1058   :   assert (rdbk == 32'h70bb2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1059   :   assert (rdbk == 32'h3615c6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1060   :   assert (rdbk == 32'h7cf932) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1061   :   assert (rdbk == 32'h7ad077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1062   :   assert (rdbk == 32'h2e013f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1063   :   assert (rdbk == 32'h76b345) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1064   :   assert (rdbk == 32'h5b5cb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1065   :   assert (rdbk == 32'h73de02) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1066   :   assert (rdbk == 32'h6389c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1067   :   assert (rdbk == 32'h4e3a95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1068   :   assert (rdbk == 32'h528dd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1069   :   assert (rdbk == 32'h22e1f9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1070   :   assert (rdbk == 32'h5fde6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1071   :   assert (rdbk == 32'h2455cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1072   :   assert (rdbk == 32'h719dc5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1073   :   assert (rdbk == 32'h4fc1e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1074   :   assert (rdbk == 32'h1ec1fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1075   :   assert (rdbk == 32'h444180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1076   :   assert (rdbk == 32'h4eaab3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1077   :   assert (rdbk == 32'h5e2e0f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1078   :   assert (rdbk == 32'h737be5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1079   :   assert (rdbk == 32'h421f37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1080   :   assert (rdbk == 32'h2a2791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1081   :   assert (rdbk == 32'h4ead5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1082   :   assert (rdbk == 32'h65216e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1083   :   assert (rdbk == 32'h38f0ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1084   :   assert (rdbk == 32'h15324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1085   :   assert (rdbk == 32'h6b23c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1086   :   assert (rdbk == 32'h3784ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1087   :   assert (rdbk == 32'h788dab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1088   :   assert (rdbk == 32'h4920ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1089   :   assert (rdbk == 32'h226677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1090   :   assert (rdbk == 32'h6fcb97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1091   :   assert (rdbk == 32'h43ce5c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1092   :   assert (rdbk == 32'h141ee8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1093   :   assert (rdbk == 32'h3a18cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1094   :   assert (rdbk == 32'h4c2578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1095   :   assert (rdbk == 32'h282bbe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1096   :   assert (rdbk == 32'h43862f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1097   :   assert (rdbk == 32'h30b57a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1098   :   assert (rdbk == 32'h1fc7b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1099   :   assert (rdbk == 32'h4f6fc2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1100   :   assert (rdbk == 32'h76489b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1101   :   assert (rdbk == 32'h4a5282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1102   :   assert (rdbk == 32'h7eba33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1103   :   assert (rdbk == 32'h1d2719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1104   :   assert (rdbk == 32'he227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1105   :   assert (rdbk == 32'h2f5739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1106   :   assert (rdbk == 32'h15472a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1107   :   assert (rdbk == 32'h5f9e51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1108   :   assert (rdbk == 32'h64aa9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1109   :   assert (rdbk == 32'h1b41d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1110   :   assert (rdbk == 32'h3145ef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1111   :   assert (rdbk == 32'h681630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1112   :   assert (rdbk == 32'h7f7546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1113   :   assert (rdbk == 32'hd4320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1114   :   assert (rdbk == 32'h2cfc92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1115   :   assert (rdbk == 32'h428dcc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1116   :   assert (rdbk == 32'h15db91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1117   :   assert (rdbk == 32'h1c476e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1118   :   assert (rdbk == 32'h48803c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1119   :   assert (rdbk == 32'h769b05) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1120   :   assert (rdbk == 32'h303fdc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1121   :   assert (rdbk == 32'h3f59f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1122   :   assert (rdbk == 32'h3ad779) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1123   :   assert (rdbk == 32'h45684c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1124   :   assert (rdbk == 32'h41e15b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1125   :   assert (rdbk == 32'h40230d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1126   :   assert (rdbk == 32'h1d6611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1127   :   assert (rdbk == 32'h626fcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1128   :   assert (rdbk == 32'h1e582c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1129   :   assert (rdbk == 32'h76bcec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1130   :   assert (rdbk == 32'h4afd27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1131   :   assert (rdbk == 32'h3c15db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1132   :   assert (rdbk == 32'h7e4efa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1133   :   assert (rdbk == 32'h2e51fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1134   :   assert (rdbk == 32'h4998ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1135   :   assert (rdbk == 32'h33f3fe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1136   :   assert (rdbk == 32'h6adc2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1137   :   assert (rdbk == 32'h51467d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1138   :   assert (rdbk == 32'h5f6808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1139   :   assert (rdbk == 32'h208d51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1140   :   assert (rdbk == 32'h30bc64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1141   :   assert (rdbk == 32'h7e76d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1142   :   assert (rdbk == 32'h3752eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1143   :   assert (rdbk == 32'h2d62be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1144   :   assert (rdbk == 32'h7a8432) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1145   :   assert (rdbk == 32'h54a4e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1146   :   assert (rdbk == 32'h12ce48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1147   :   assert (rdbk == 32'h34dad6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1148   :   assert (rdbk == 32'h7d8204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1149   :   assert (rdbk == 32'h49b2f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1150   :   assert (rdbk == 32'h1bb9e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1151   :   assert (rdbk == 32'h243eb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1152   :   assert (rdbk == 32'h666a5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1153   :   assert (rdbk == 32'h15de00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1154   :   assert (rdbk == 32'h668189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1155   :   assert (rdbk == 32'h386878) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1156   :   assert (rdbk == 32'h1941d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1157   :   assert (rdbk == 32'h162447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1158   :   assert (rdbk == 32'h5d4c39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1159   :   assert (rdbk == 32'h4f7a30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1160   :   assert (rdbk == 32'h69834c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1161   :   assert (rdbk == 32'h4e44b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1162   :   assert (rdbk == 32'h6c2e0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1163   :   assert (rdbk == 32'h674ac8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1164   :   assert (rdbk == 32'h388bea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1165   :   assert (rdbk == 32'h7f6c12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1166   :   assert (rdbk == 32'h235752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1167   :   assert (rdbk == 32'h32c1f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1168   :   assert (rdbk == 32'h7a54cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1169   :   assert (rdbk == 32'h446124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1170   :   assert (rdbk == 32'h4995b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1171   :   assert (rdbk == 32'h315386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1172   :   assert (rdbk == 32'h583f07) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1173   :   assert (rdbk == 32'h78e84b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1174   :   assert (rdbk == 32'h7a4629) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1175   :   assert (rdbk == 32'h78dee9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1176   :   assert (rdbk == 32'h4b7602) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1177   :   assert (rdbk == 32'h25c289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1178   :   assert (rdbk == 32'h54c59e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1179   :   assert (rdbk == 32'h640020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1180   :   assert (rdbk == 32'h5b94d9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1181   :   assert (rdbk == 32'h39474c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1182   :   assert (rdbk == 32'h7f3c56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1183   :   assert (rdbk == 32'h62dd2a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1184   :   assert (rdbk == 32'h51b0f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1185   :   assert (rdbk == 32'h36aa31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1186   :   assert (rdbk == 32'h3beed8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1187   :   assert (rdbk == 32'h1d4f9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1188   :   assert (rdbk == 32'h70a664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1189   :   assert (rdbk == 32'h297a4e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1190   :   assert (rdbk == 32'h4fcb87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1191   :   assert (rdbk == 32'ha129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1192   :   assert (rdbk == 32'h9e709) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1193   :   assert (rdbk == 32'ha4cc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1194   :   assert (rdbk == 32'h1e0574) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1195   :   assert (rdbk == 32'h3b8334) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1196   :   assert (rdbk == 32'h72f174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1197   :   assert (rdbk == 32'h58e433) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1198   :   assert (rdbk == 32'h41196d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1199   :   assert (rdbk == 32'h6751c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1200   :   assert (rdbk == 32'h11a0ae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1201   :   assert (rdbk == 32'h224223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1202   :   assert (rdbk == 32'h754e0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1203   :   assert (rdbk == 32'h233922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1204   :   assert (rdbk == 32'h7b6ffb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1205   :   assert (rdbk == 32'h855e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1206   :   assert (rdbk == 32'h2502fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1207   :   assert (rdbk == 32'h2931c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1208   :   assert (rdbk == 32'h2a55de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1209   :   assert (rdbk == 32'h22a30d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1210   :   assert (rdbk == 32'h93cce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1211   :   assert (rdbk == 32'h4fd2f8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1212   :   assert (rdbk == 32'h36a4cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1213   :   assert (rdbk == 32'h40d574) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1214   :   assert (rdbk == 32'h1d873d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1215   :   assert (rdbk == 32'h5b227f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1216   :   assert (rdbk == 32'h6c7b15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1217   :   assert (rdbk == 32'h48a6c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1218   :   assert (rdbk == 32'h491ded) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1219   :   assert (rdbk == 32'h5a87c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1220   :   assert (rdbk == 32'h24c105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1221   :   assert (rdbk == 32'h3417d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1222   :   assert (rdbk == 32'h69c9fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1223   :   assert (rdbk == 32'h5525b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1224   :   assert (rdbk == 32'h64ff24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1225   :   assert (rdbk == 32'h567a90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1226   :   assert (rdbk == 32'h381a0f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1227   :   assert (rdbk == 32'h4c602a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1228   :   assert (rdbk == 32'h53e6ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1229   :   assert (rdbk == 32'h7ea2db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1230   :   assert (rdbk == 32'h6ed52c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1231   :   assert (rdbk == 32'h11553f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1232   :   assert (rdbk == 32'h18f4db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1233   :   assert (rdbk == 32'h5b172f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1234   :   assert (rdbk == 32'h1f8138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1235   :   assert (rdbk == 32'h3e7b8d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1236   :   assert (rdbk == 32'h70ff94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1237   :   assert (rdbk == 32'h59beaf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1238   :   assert (rdbk == 32'h2736a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1239   :   assert (rdbk == 32'h630633) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1240   :   assert (rdbk == 32'h16bfcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1241   :   assert (rdbk == 32'h76ff0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1242   :   assert (rdbk == 32'h7e7b28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1243   :   assert (rdbk == 32'h5a30a1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1244   :   assert (rdbk == 32'h3c584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1245   :   assert (rdbk == 32'h2e4843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1246   :   assert (rdbk == 32'h3c483e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1247   :   assert (rdbk == 32'h2289d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1248   :   assert (rdbk == 32'h4e9ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1249   :   assert (rdbk == 32'h4ddc23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1250   :   assert (rdbk == 32'h3b01da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1251   :   assert (rdbk == 32'h11086b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1252   :   assert (rdbk == 32'h16eb1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1253   :   assert (rdbk == 32'h30f4f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1254   :   assert (rdbk == 32'h33e0bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1255   :   assert (rdbk == 32'h635165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1256   :   assert (rdbk == 32'h335f22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1257   :   assert (rdbk == 32'h6559a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1258   :   assert (rdbk == 32'h72eb9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1259   :   assert (rdbk == 32'h5b4907) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1260   :   assert (rdbk == 32'h6a44a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1261   :   assert (rdbk == 32'h1847aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1262   :   assert (rdbk == 32'h4c072a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1263   :   assert (rdbk == 32'h2ae0e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1264   :   assert (rdbk == 32'hd385f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1265   :   assert (rdbk == 32'h2e3f2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1266   :   assert (rdbk == 32'h5bdbaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1267   :   assert (rdbk == 32'h1b5438) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1268   :   assert (rdbk == 32'h563d07) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1269   :   assert (rdbk == 32'hfb2df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1270   :   assert (rdbk == 32'h4073a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1271   :   assert (rdbk == 32'h3f8b46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1272   :   assert (rdbk == 32'h534a1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1273   :   assert (rdbk == 32'h50047e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1274   :   assert (rdbk == 32'h184c8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1275   :   assert (rdbk == 32'h5fc6ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1276   :   assert (rdbk == 32'h4f0e58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1277   :   assert (rdbk == 32'h271052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1278   :   assert (rdbk == 32'h5eb4d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1279   :   assert (rdbk == 32'h4cfe50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h101
	1280   :   assert (rdbk == 32'h6fe933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1281   :   assert (rdbk == 32'h6b3ff4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1282   :   assert (rdbk == 32'h51bd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1283   :   assert (rdbk == 32'h3e0a60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1284   :   assert (rdbk == 32'h58a83b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1285   :   assert (rdbk == 32'h2170ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1286   :   assert (rdbk == 32'h3c8137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1287   :   assert (rdbk == 32'h32b38c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1288   :   assert (rdbk == 32'h5654f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1289   :   assert (rdbk == 32'h63a1b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1290   :   assert (rdbk == 32'h49cc3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1291   :   assert (rdbk == 32'h23cd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1292   :   assert (rdbk == 32'h6f3767) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1293   :   assert (rdbk == 32'h3932ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1294   :   assert (rdbk == 32'h25a89e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1295   :   assert (rdbk == 32'h79d98c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1296   :   assert (rdbk == 32'he75d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1297   :   assert (rdbk == 32'h33fe18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1298   :   assert (rdbk == 32'h36339e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1299   :   assert (rdbk == 32'h58e8da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1300   :   assert (rdbk == 32'h7e97ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1301   :   assert (rdbk == 32'h12d506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1302   :   assert (rdbk == 32'h75a18b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1303   :   assert (rdbk == 32'h1eda70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1304   :   assert (rdbk == 32'h18c0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1305   :   assert (rdbk == 32'h78083f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1306   :   assert (rdbk == 32'h372b91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1307   :   assert (rdbk == 32'h2917ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1308   :   assert (rdbk == 32'h345e96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1309   :   assert (rdbk == 32'h15ed56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1310   :   assert (rdbk == 32'h2cea63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1311   :   assert (rdbk == 32'h577536) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1312   :   assert (rdbk == 32'h74df5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1313   :   assert (rdbk == 32'h446c5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1314   :   assert (rdbk == 32'h2c829c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1315   :   assert (rdbk == 32'h5fee74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1316   :   assert (rdbk == 32'h1a5bb0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1317   :   assert (rdbk == 32'h431eee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1318   :   assert (rdbk == 32'h61eb0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1319   :   assert (rdbk == 32'h262405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1320   :   assert (rdbk == 32'h2781f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1321   :   assert (rdbk == 32'h667f58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1322   :   assert (rdbk == 32'h544f7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1323   :   assert (rdbk == 32'h138728) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1324   :   assert (rdbk == 32'h55ad45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1325   :   assert (rdbk == 32'h697ec9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1326   :   assert (rdbk == 32'h27caf7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1327   :   assert (rdbk == 32'h4e4108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1328   :   assert (rdbk == 32'hc7bda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1329   :   assert (rdbk == 32'h147bb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1330   :   assert (rdbk == 32'h10a4b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1331   :   assert (rdbk == 32'h42beca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1332   :   assert (rdbk == 32'he1b63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1333   :   assert (rdbk == 32'hf3ea9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1334   :   assert (rdbk == 32'h67b147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1335   :   assert (rdbk == 32'h3ec3dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1336   :   assert (rdbk == 32'h7d9be3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1337   :   assert (rdbk == 32'h4211e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1338   :   assert (rdbk == 32'h55a463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1339   :   assert (rdbk == 32'h6f4a84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1340   :   assert (rdbk == 32'h6cf8a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1341   :   assert (rdbk == 32'h5feb21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1342   :   assert (rdbk == 32'h52685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1343   :   assert (rdbk == 32'h7350f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1344   :   assert (rdbk == 32'h474b1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1345   :   assert (rdbk == 32'h396a58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1346   :   assert (rdbk == 32'h182c87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1347   :   assert (rdbk == 32'h1aa6ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1348   :   assert (rdbk == 32'h3771c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1349   :   assert (rdbk == 32'h7b1256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1350   :   assert (rdbk == 32'h752f6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1351   :   assert (rdbk == 32'h482a5e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1352   :   assert (rdbk == 32'h6ac466) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1353   :   assert (rdbk == 32'h42b700) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1354   :   assert (rdbk == 32'h59f440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1355   :   assert (rdbk == 32'h33d193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1356   :   assert (rdbk == 32'h64a842) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1357   :   assert (rdbk == 32'h5161ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1358   :   assert (rdbk == 32'h25a521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1359   :   assert (rdbk == 32'h4bb894) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1360   :   assert (rdbk == 32'h7a5e60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1361   :   assert (rdbk == 32'h62a488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1362   :   assert (rdbk == 32'h680ce5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1363   :   assert (rdbk == 32'h57cdbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1364   :   assert (rdbk == 32'h53e9f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1365   :   assert (rdbk == 32'h64d2d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1366   :   assert (rdbk == 32'h739bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1367   :   assert (rdbk == 32'h7a1af1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1368   :   assert (rdbk == 32'h4b7d8e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1369   :   assert (rdbk == 32'h6a0ea5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1370   :   assert (rdbk == 32'h389c56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1371   :   assert (rdbk == 32'h285c36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1372   :   assert (rdbk == 32'h36ee92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1373   :   assert (rdbk == 32'h2b5d0f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1374   :   assert (rdbk == 32'h54a07d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1375   :   assert (rdbk == 32'h16816e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1376   :   assert (rdbk == 32'h30e5a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1377   :   assert (rdbk == 32'h1796ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1378   :   assert (rdbk == 32'h1c38fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1379   :   assert (rdbk == 32'h64adb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1380   :   assert (rdbk == 32'h24bc58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1381   :   assert (rdbk == 32'h4cb5fe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1382   :   assert (rdbk == 32'h4e2ef9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1383   :   assert (rdbk == 32'h7c00ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1384   :   assert (rdbk == 32'h33fa54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1385   :   assert (rdbk == 32'h475c26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1386   :   assert (rdbk == 32'h76ae92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1387   :   assert (rdbk == 32'h33365c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1388   :   assert (rdbk == 32'h1b832f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1389   :   assert (rdbk == 32'h6c0867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1390   :   assert (rdbk == 32'h27b0ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1391   :   assert (rdbk == 32'h5136d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1392   :   assert (rdbk == 32'h4d536e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1393   :   assert (rdbk == 32'h7cb2a4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1394   :   assert (rdbk == 32'h4b3d59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1395   :   assert (rdbk == 32'h3e0e95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1396   :   assert (rdbk == 32'h47db34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1397   :   assert (rdbk == 32'h4eb5b2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1398   :   assert (rdbk == 32'h33c032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1399   :   assert (rdbk == 32'h769e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1400   :   assert (rdbk == 32'hfba9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1401   :   assert (rdbk == 32'h4e462b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1402   :   assert (rdbk == 32'h11eef6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1403   :   assert (rdbk == 32'h4cf583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1404   :   assert (rdbk == 32'h505212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1405   :   assert (rdbk == 32'h1736a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1406   :   assert (rdbk == 32'h6f3bb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1407   :   assert (rdbk == 32'h6405bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1408   :   assert (rdbk == 32'h6ff6a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1409   :   assert (rdbk == 32'h4d104f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1410   :   assert (rdbk == 32'h11de5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1411   :   assert (rdbk == 32'h333f67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1412   :   assert (rdbk == 32'hf3286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1413   :   assert (rdbk == 32'h6dee15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1414   :   assert (rdbk == 32'h36f8cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1415   :   assert (rdbk == 32'h71de6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1416   :   assert (rdbk == 32'h4ac94e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1417   :   assert (rdbk == 32'h5a0ff3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1418   :   assert (rdbk == 32'h2a1a88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1419   :   assert (rdbk == 32'h183b75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1420   :   assert (rdbk == 32'h67ebe7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1421   :   assert (rdbk == 32'h5c2d24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1422   :   assert (rdbk == 32'h519be1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1423   :   assert (rdbk == 32'h5c12c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1424   :   assert (rdbk == 32'h3b50b2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1425   :   assert (rdbk == 32'h117476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1426   :   assert (rdbk == 32'h146965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1427   :   assert (rdbk == 32'h48f8dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1428   :   assert (rdbk == 32'h62fe27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1429   :   assert (rdbk == 32'h7cf6de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1430   :   assert (rdbk == 32'h75fcad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1431   :   assert (rdbk == 32'hce8d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1432   :   assert (rdbk == 32'h213bab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1433   :   assert (rdbk == 32'h17c95c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1434   :   assert (rdbk == 32'h5d8ee0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1435   :   assert (rdbk == 32'h552a15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1436   :   assert (rdbk == 32'h7f4477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1437   :   assert (rdbk == 32'h2f39aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1438   :   assert (rdbk == 32'h60dc7b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1439   :   assert (rdbk == 32'h5d0b43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1440   :   assert (rdbk == 32'hed1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1441   :   assert (rdbk == 32'h53eb42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1442   :   assert (rdbk == 32'hc287b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1443   :   assert (rdbk == 32'h23d91f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1444   :   assert (rdbk == 32'h530605) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1445   :   assert (rdbk == 32'h421bcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1446   :   assert (rdbk == 32'h596ffb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1447   :   assert (rdbk == 32'hdb517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1448   :   assert (rdbk == 32'hff10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1449   :   assert (rdbk == 32'h508399) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1450   :   assert (rdbk == 32'h387e7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1451   :   assert (rdbk == 32'h9caa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1452   :   assert (rdbk == 32'h41cca8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1453   :   assert (rdbk == 32'h50e6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1454   :   assert (rdbk == 32'h4d213a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1455   :   assert (rdbk == 32'h10c609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1456   :   assert (rdbk == 32'h617eff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1457   :   assert (rdbk == 32'h4de692) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1458   :   assert (rdbk == 32'h1c0dea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1459   :   assert (rdbk == 32'h4a7253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1460   :   assert (rdbk == 32'h696924) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1461   :   assert (rdbk == 32'h4c2686) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1462   :   assert (rdbk == 32'h6297c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1463   :   assert (rdbk == 32'h74ed9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1464   :   assert (rdbk == 32'h4437c6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1465   :   assert (rdbk == 32'h6b156a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1466   :   assert (rdbk == 32'h34209e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1467   :   assert (rdbk == 32'h26d8bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1468   :   assert (rdbk == 32'h4f86c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1469   :   assert (rdbk == 32'h40eaf6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1470   :   assert (rdbk == 32'hc672b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1471   :   assert (rdbk == 32'h3aa6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1472   :   assert (rdbk == 32'h13b826) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1473   :   assert (rdbk == 32'h4e4299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1474   :   assert (rdbk == 32'h2389e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1475   :   assert (rdbk == 32'h23bb8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1476   :   assert (rdbk == 32'h7d08de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1477   :   assert (rdbk == 32'h5b54e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1478   :   assert (rdbk == 32'h78f686) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1479   :   assert (rdbk == 32'h25d73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1480   :   assert (rdbk == 32'h1304eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1481   :   assert (rdbk == 32'h4178b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1482   :   assert (rdbk == 32'h751660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1483   :   assert (rdbk == 32'h774a58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1484   :   assert (rdbk == 32'h1d967) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1485   :   assert (rdbk == 32'h78059d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1486   :   assert (rdbk == 32'h6ffbd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1487   :   assert (rdbk == 32'h530241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1488   :   assert (rdbk == 32'h21b06) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1489   :   assert (rdbk == 32'h59dac4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1490   :   assert (rdbk == 32'h3c4e04) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1491   :   assert (rdbk == 32'h573588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1492   :   assert (rdbk == 32'h249954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1493   :   assert (rdbk == 32'h75c9b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1494   :   assert (rdbk == 32'h2bb577) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1495   :   assert (rdbk == 32'h35416a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1496   :   assert (rdbk == 32'h64faaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1497   :   assert (rdbk == 32'h37b4ef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1498   :   assert (rdbk == 32'h200694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1499   :   assert (rdbk == 32'h5c0309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1500   :   assert (rdbk == 32'h2ada76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1501   :   assert (rdbk == 32'h48a144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1502   :   assert (rdbk == 32'h5b8215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1503   :   assert (rdbk == 32'hc044b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1504   :   assert (rdbk == 32'h5e446f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1505   :   assert (rdbk == 32'h33d78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1506   :   assert (rdbk == 32'hda812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1507   :   assert (rdbk == 32'h3b44c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1508   :   assert (rdbk == 32'h760f09) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1509   :   assert (rdbk == 32'h87944) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1510   :   assert (rdbk == 32'h3bdc3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1511   :   assert (rdbk == 32'h4d7b5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1512   :   assert (rdbk == 32'h705a60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1513   :   assert (rdbk == 32'h60ec3b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1514   :   assert (rdbk == 32'he2413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1515   :   assert (rdbk == 32'h2a513f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1516   :   assert (rdbk == 32'h203288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1517   :   assert (rdbk == 32'h6ae4fe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1518   :   assert (rdbk == 32'h140722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1519   :   assert (rdbk == 32'h706086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1520   :   assert (rdbk == 32'h1c5982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1521   :   assert (rdbk == 32'h71b666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1522   :   assert (rdbk == 32'h73521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1523   :   assert (rdbk == 32'hefd13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1524   :   assert (rdbk == 32'h423384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1525   :   assert (rdbk == 32'h42f12f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1526   :   assert (rdbk == 32'h2e5516) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1527   :   assert (rdbk == 32'h1344bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1528   :   assert (rdbk == 32'h4d11ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1529   :   assert (rdbk == 32'h5383f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1530   :   assert (rdbk == 32'h3c5d95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1531   :   assert (rdbk == 32'h2571c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1532   :   assert (rdbk == 32'h2a3144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1533   :   assert (rdbk == 32'h122ce4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1534   :   assert (rdbk == 32'h747023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1535   :   assert (rdbk == 32'h6e77fe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h102
	1536   :   assert (rdbk == 32'h692c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1537   :   assert (rdbk == 32'h278b92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1538   :   assert (rdbk == 32'h16563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1539   :   assert (rdbk == 32'h1da7f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1540   :   assert (rdbk == 32'h23a853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1541   :   assert (rdbk == 32'hc3c72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1542   :   assert (rdbk == 32'h3b0c63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1543   :   assert (rdbk == 32'h180e79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1544   :   assert (rdbk == 32'h7666b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1545   :   assert (rdbk == 32'h1b7dc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1546   :   assert (rdbk == 32'h445de8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1547   :   assert (rdbk == 32'h1faa50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1548   :   assert (rdbk == 32'h51aac7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1549   :   assert (rdbk == 32'h59eed4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1550   :   assert (rdbk == 32'h40dbe4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1551   :   assert (rdbk == 32'h1d69f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1552   :   assert (rdbk == 32'h76fe9e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1553   :   assert (rdbk == 32'h27be06) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1554   :   assert (rdbk == 32'hfd9aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1555   :   assert (rdbk == 32'h4aafcd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1556   :   assert (rdbk == 32'h29fdf9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1557   :   assert (rdbk == 32'h48cdf8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1558   :   assert (rdbk == 32'hf01af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1559   :   assert (rdbk == 32'h2de771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1560   :   assert (rdbk == 32'h4ebe75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1561   :   assert (rdbk == 32'h308d79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1562   :   assert (rdbk == 32'h3a56b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1563   :   assert (rdbk == 32'h76eb3e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1564   :   assert (rdbk == 32'h371136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1565   :   assert (rdbk == 32'h38c919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1566   :   assert (rdbk == 32'he6cee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1567   :   assert (rdbk == 32'h4043c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1568   :   assert (rdbk == 32'h1b57f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1569   :   assert (rdbk == 32'h554d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1570   :   assert (rdbk == 32'h26a9eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1571   :   assert (rdbk == 32'h15d900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1572   :   assert (rdbk == 32'h3f0a26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1573   :   assert (rdbk == 32'h42f22b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1574   :   assert (rdbk == 32'h7ba94e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1575   :   assert (rdbk == 32'h36709b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1576   :   assert (rdbk == 32'h14891e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1577   :   assert (rdbk == 32'h31bd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1578   :   assert (rdbk == 32'h1d09e2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1579   :   assert (rdbk == 32'h1eb3ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1580   :   assert (rdbk == 32'h2a6af7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1581   :   assert (rdbk == 32'h7885e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1582   :   assert (rdbk == 32'h5e4892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1583   :   assert (rdbk == 32'h4ec435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1584   :   assert (rdbk == 32'h5eb9e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1585   :   assert (rdbk == 32'h4dfbda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1586   :   assert (rdbk == 32'h6e77f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1587   :   assert (rdbk == 32'h23a02f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1588   :   assert (rdbk == 32'h131306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1589   :   assert (rdbk == 32'h659a14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1590   :   assert (rdbk == 32'h7d4677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1591   :   assert (rdbk == 32'h63530c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1592   :   assert (rdbk == 32'h16d2bf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1593   :   assert (rdbk == 32'h2c54d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1594   :   assert (rdbk == 32'h3f1015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1595   :   assert (rdbk == 32'h126365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1596   :   assert (rdbk == 32'h5d6e11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1597   :   assert (rdbk == 32'h182d1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1598   :   assert (rdbk == 32'h5b343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1599   :   assert (rdbk == 32'h347dec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1600   :   assert (rdbk == 32'h1903a4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1601   :   assert (rdbk == 32'h320fc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1602   :   assert (rdbk == 32'h64abbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1603   :   assert (rdbk == 32'h470813) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1604   :   assert (rdbk == 32'h5d586f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1605   :   assert (rdbk == 32'h6ead88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1606   :   assert (rdbk == 32'h6070ef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1607   :   assert (rdbk == 32'h30210c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1608   :   assert (rdbk == 32'h394b59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1609   :   assert (rdbk == 32'h48050b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1610   :   assert (rdbk == 32'h38a8e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1611   :   assert (rdbk == 32'h1d79fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1612   :   assert (rdbk == 32'h2c1ff6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1613   :   assert (rdbk == 32'h7e78ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1614   :   assert (rdbk == 32'h14fba9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1615   :   assert (rdbk == 32'h3f6e86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1616   :   assert (rdbk == 32'h15eafe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1617   :   assert (rdbk == 32'h365c25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1618   :   assert (rdbk == 32'h563e0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1619   :   assert (rdbk == 32'h79ecaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1620   :   assert (rdbk == 32'h264f9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1621   :   assert (rdbk == 32'h71e5c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1622   :   assert (rdbk == 32'h77ecb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1623   :   assert (rdbk == 32'h69cc30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1624   :   assert (rdbk == 32'h68c8bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1625   :   assert (rdbk == 32'h177e1e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1626   :   assert (rdbk == 32'h733845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1627   :   assert (rdbk == 32'h6465cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1628   :   assert (rdbk == 32'h6ecbd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1629   :   assert (rdbk == 32'h2c0c72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1630   :   assert (rdbk == 32'h1fdaa5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1631   :   assert (rdbk == 32'hffb89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1632   :   assert (rdbk == 32'h7e5aa7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1633   :   assert (rdbk == 32'h36b898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1634   :   assert (rdbk == 32'h7081b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1635   :   assert (rdbk == 32'h24b0ec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1636   :   assert (rdbk == 32'h32053) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1637   :   assert (rdbk == 32'h515dfb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1638   :   assert (rdbk == 32'h7c1c58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1639   :   assert (rdbk == 32'h74e6c4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1640   :   assert (rdbk == 32'h75c840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1641   :   assert (rdbk == 32'h3de4ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1642   :   assert (rdbk == 32'hff953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1643   :   assert (rdbk == 32'h188de0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1644   :   assert (rdbk == 32'h6b55f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1645   :   assert (rdbk == 32'h1a19ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1646   :   assert (rdbk == 32'h90a3e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1647   :   assert (rdbk == 32'h33b009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1648   :   assert (rdbk == 32'h28cef1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1649   :   assert (rdbk == 32'h274b18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1650   :   assert (rdbk == 32'h43e284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1651   :   assert (rdbk == 32'h4bb893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1652   :   assert (rdbk == 32'h3c944d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1653   :   assert (rdbk == 32'h36a30d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1654   :   assert (rdbk == 32'h655fd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1655   :   assert (rdbk == 32'h7b9a1a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1656   :   assert (rdbk == 32'h412d82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1657   :   assert (rdbk == 32'h72703c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1658   :   assert (rdbk == 32'h68a15f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1659   :   assert (rdbk == 32'h380849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1660   :   assert (rdbk == 32'h5dea24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1661   :   assert (rdbk == 32'h24de06) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1662   :   assert (rdbk == 32'h2200b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1663   :   assert (rdbk == 32'h4bbe14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1664   :   assert (rdbk == 32'h2f6008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1665   :   assert (rdbk == 32'hc6b6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1666   :   assert (rdbk == 32'h7ec2e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1667   :   assert (rdbk == 32'h5e1b2b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1668   :   assert (rdbk == 32'h112e4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1669   :   assert (rdbk == 32'h66ecb7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1670   :   assert (rdbk == 32'h796a69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1671   :   assert (rdbk == 32'h75bf19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1672   :   assert (rdbk == 32'h793633) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1673   :   assert (rdbk == 32'h3850ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1674   :   assert (rdbk == 32'h2f340) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1675   :   assert (rdbk == 32'h412f46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1676   :   assert (rdbk == 32'h62de3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1677   :   assert (rdbk == 32'h60ccf4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1678   :   assert (rdbk == 32'h49fd30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1679   :   assert (rdbk == 32'h168db8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1680   :   assert (rdbk == 32'h92c63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1681   :   assert (rdbk == 32'h22fde7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1682   :   assert (rdbk == 32'hdbd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1683   :   assert (rdbk == 32'h2fbff3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1684   :   assert (rdbk == 32'h3eb70c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1685   :   assert (rdbk == 32'h285e86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1686   :   assert (rdbk == 32'h39355a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1687   :   assert (rdbk == 32'h62cb95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1688   :   assert (rdbk == 32'h29e4a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1689   :   assert (rdbk == 32'h57deef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1690   :   assert (rdbk == 32'h57d88e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1691   :   assert (rdbk == 32'h1298d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1692   :   assert (rdbk == 32'h6d4860) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1693   :   assert (rdbk == 32'h605faf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1694   :   assert (rdbk == 32'h637b00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1695   :   assert (rdbk == 32'h2a28d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1696   :   assert (rdbk == 32'h2d9771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1697   :   assert (rdbk == 32'h2d30f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1698   :   assert (rdbk == 32'hffe30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1699   :   assert (rdbk == 32'h6a6b1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1700   :   assert (rdbk == 32'h5f5903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1701   :   assert (rdbk == 32'h5f3c11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1702   :   assert (rdbk == 32'h4ca7be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1703   :   assert (rdbk == 32'h5d5bb0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1704   :   assert (rdbk == 32'h2b12b1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1705   :   assert (rdbk == 32'h5f46d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1706   :   assert (rdbk == 32'h7383d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1707   :   assert (rdbk == 32'h6e48a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1708   :   assert (rdbk == 32'h24be69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1709   :   assert (rdbk == 32'h2ca36a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1710   :   assert (rdbk == 32'h2d5ee2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1711   :   assert (rdbk == 32'h15c8f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1712   :   assert (rdbk == 32'h5cda7c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1713   :   assert (rdbk == 32'h339f56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1714   :   assert (rdbk == 32'h60b0be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1715   :   assert (rdbk == 32'h3b01de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1716   :   assert (rdbk == 32'h636071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1717   :   assert (rdbk == 32'h2822de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1718   :   assert (rdbk == 32'h6108f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1719   :   assert (rdbk == 32'h7e2405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1720   :   assert (rdbk == 32'h71ad06) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1721   :   assert (rdbk == 32'h5b323e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1722   :   assert (rdbk == 32'h645880) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1723   :   assert (rdbk == 32'h3ea7ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1724   :   assert (rdbk == 32'h5c34a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1725   :   assert (rdbk == 32'h25765c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1726   :   assert (rdbk == 32'h32e6f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1727   :   assert (rdbk == 32'h5a0c61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1728   :   assert (rdbk == 32'h41acb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1729   :   assert (rdbk == 32'h6afd3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1730   :   assert (rdbk == 32'h51c0eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1731   :   assert (rdbk == 32'h333d76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1732   :   assert (rdbk == 32'h4986c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1733   :   assert (rdbk == 32'h305479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1734   :   assert (rdbk == 32'h4dfd7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1735   :   assert (rdbk == 32'h7a6fda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1736   :   assert (rdbk == 32'h2342ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1737   :   assert (rdbk == 32'h58a6c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1738   :   assert (rdbk == 32'h6e6b6b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1739   :   assert (rdbk == 32'h4831ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1740   :   assert (rdbk == 32'h50721e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1741   :   assert (rdbk == 32'h710321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1742   :   assert (rdbk == 32'h645242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1743   :   assert (rdbk == 32'hcbc84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1744   :   assert (rdbk == 32'h3d939c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1745   :   assert (rdbk == 32'h5b99be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1746   :   assert (rdbk == 32'h44f004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1747   :   assert (rdbk == 32'h1f9cdb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1748   :   assert (rdbk == 32'h650920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1749   :   assert (rdbk == 32'h376b55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1750   :   assert (rdbk == 32'h3a2399) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1751   :   assert (rdbk == 32'h771f1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1752   :   assert (rdbk == 32'hececc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1753   :   assert (rdbk == 32'h34435e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1754   :   assert (rdbk == 32'h73efdb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1755   :   assert (rdbk == 32'h77fcb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1756   :   assert (rdbk == 32'h46c91f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1757   :   assert (rdbk == 32'h7b993e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1758   :   assert (rdbk == 32'h2a18df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1759   :   assert (rdbk == 32'h5d552b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1760   :   assert (rdbk == 32'h2662d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1761   :   assert (rdbk == 32'h1b2923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1762   :   assert (rdbk == 32'h340f18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1763   :   assert (rdbk == 32'h2a6e19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1764   :   assert (rdbk == 32'h709540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1765   :   assert (rdbk == 32'h86a5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1766   :   assert (rdbk == 32'h483b33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1767   :   assert (rdbk == 32'h34f00f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1768   :   assert (rdbk == 32'h77bc99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1769   :   assert (rdbk == 32'h2864d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1770   :   assert (rdbk == 32'h51590c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1771   :   assert (rdbk == 32'h18bf50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1772   :   assert (rdbk == 32'h9dbd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1773   :   assert (rdbk == 32'hd9ddf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1774   :   assert (rdbk == 32'h319d87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1775   :   assert (rdbk == 32'h1028d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1776   :   assert (rdbk == 32'h43d73e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1777   :   assert (rdbk == 32'h6fa300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1778   :   assert (rdbk == 32'h19d9d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1779   :   assert (rdbk == 32'h239272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1780   :   assert (rdbk == 32'h12c204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1781   :   assert (rdbk == 32'h508bbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1782   :   assert (rdbk == 32'h40d2c4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1783   :   assert (rdbk == 32'h527bfd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1784   :   assert (rdbk == 32'h3221a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1785   :   assert (rdbk == 32'h3a4ce4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1786   :   assert (rdbk == 32'h49e290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1787   :   assert (rdbk == 32'h55eb8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1788   :   assert (rdbk == 32'h655b55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1789   :   assert (rdbk == 32'h220d45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1790   :   assert (rdbk == 32'h54d758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1791   :   assert (rdbk == 32'h370594) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h103
	1792   :   assert (rdbk == 32'h4ce166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1793   :   assert (rdbk == 32'h61ea71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1794   :   assert (rdbk == 32'he3e8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1795   :   assert (rdbk == 32'h69e393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1796   :   assert (rdbk == 32'h65ccea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1797   :   assert (rdbk == 32'h36baa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1798   :   assert (rdbk == 32'h71b9d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1799   :   assert (rdbk == 32'h309e01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1800   :   assert (rdbk == 32'h1c1c7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1801   :   assert (rdbk == 32'h5e17c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1802   :   assert (rdbk == 32'h47035a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1803   :   assert (rdbk == 32'h456087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1804   :   assert (rdbk == 32'hdf6ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1805   :   assert (rdbk == 32'h55ffd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1806   :   assert (rdbk == 32'h222eca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1807   :   assert (rdbk == 32'hba26f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1808   :   assert (rdbk == 32'h161818) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1809   :   assert (rdbk == 32'h2315d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1810   :   assert (rdbk == 32'h1bd399) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1811   :   assert (rdbk == 32'h35450f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1812   :   assert (rdbk == 32'h7dbde7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1813   :   assert (rdbk == 32'h3b2d52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1814   :   assert (rdbk == 32'h3135fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1815   :   assert (rdbk == 32'hbbcf3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1816   :   assert (rdbk == 32'h7c0b70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1817   :   assert (rdbk == 32'h66387e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1818   :   assert (rdbk == 32'h4ff71f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1819   :   assert (rdbk == 32'h223f4d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1820   :   assert (rdbk == 32'he1ed5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1821   :   assert (rdbk == 32'h271fa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1822   :   assert (rdbk == 32'hc9a54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1823   :   assert (rdbk == 32'h560f00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1824   :   assert (rdbk == 32'h39d2a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1825   :   assert (rdbk == 32'h1504be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1826   :   assert (rdbk == 32'h2cdad9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1827   :   assert (rdbk == 32'h28cab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1828   :   assert (rdbk == 32'h643003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1829   :   assert (rdbk == 32'h5b2862) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1830   :   assert (rdbk == 32'h463f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1831   :   assert (rdbk == 32'h7f2c78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1832   :   assert (rdbk == 32'h7054da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1833   :   assert (rdbk == 32'h1cb81d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1834   :   assert (rdbk == 32'h1a2408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1835   :   assert (rdbk == 32'h4123a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1836   :   assert (rdbk == 32'h5d88b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1837   :   assert (rdbk == 32'h3b9d8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1838   :   assert (rdbk == 32'h2793bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1839   :   assert (rdbk == 32'h1b1a5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1840   :   assert (rdbk == 32'h6fb818) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1841   :   assert (rdbk == 32'h338873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1842   :   assert (rdbk == 32'h78eb5c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1843   :   assert (rdbk == 32'h609fce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1844   :   assert (rdbk == 32'h3c7f7a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1845   :   assert (rdbk == 32'h2e6b4c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1846   :   assert (rdbk == 32'h273c81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1847   :   assert (rdbk == 32'h30e8a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1848   :   assert (rdbk == 32'h730b2f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1849   :   assert (rdbk == 32'h6543ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1850   :   assert (rdbk == 32'h2da46b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1851   :   assert (rdbk == 32'h595cd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1852   :   assert (rdbk == 32'h7db795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1853   :   assert (rdbk == 32'h131c6b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1854   :   assert (rdbk == 32'h713b87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1855   :   assert (rdbk == 32'h44ee14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1856   :   assert (rdbk == 32'hc47b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1857   :   assert (rdbk == 32'h2d6264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1858   :   assert (rdbk == 32'h4ec349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1859   :   assert (rdbk == 32'h3d5998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1860   :   assert (rdbk == 32'h22afc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1861   :   assert (rdbk == 32'h4beef2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1862   :   assert (rdbk == 32'h50466e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1863   :   assert (rdbk == 32'h67beb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1864   :   assert (rdbk == 32'h208f0f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1865   :   assert (rdbk == 32'h4ed8fe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1866   :   assert (rdbk == 32'h3cf08c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1867   :   assert (rdbk == 32'h6deb08) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1868   :   assert (rdbk == 32'h223c78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1869   :   assert (rdbk == 32'h4e1579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1870   :   assert (rdbk == 32'hc0706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1871   :   assert (rdbk == 32'h66491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1872   :   assert (rdbk == 32'h31ab17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1873   :   assert (rdbk == 32'h4995e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1874   :   assert (rdbk == 32'h3a295f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1875   :   assert (rdbk == 32'h3d5f73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1876   :   assert (rdbk == 32'h474d4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1877   :   assert (rdbk == 32'h289b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1878   :   assert (rdbk == 32'h57d9fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1879   :   assert (rdbk == 32'h1b9b59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1880   :   assert (rdbk == 32'h49ed87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1881   :   assert (rdbk == 32'h767914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1882   :   assert (rdbk == 32'h4966db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1883   :   assert (rdbk == 32'h1b1316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1884   :   assert (rdbk == 32'h2e60f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1885   :   assert (rdbk == 32'h2c035e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1886   :   assert (rdbk == 32'h72e2a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1887   :   assert (rdbk == 32'h63c54c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1888   :   assert (rdbk == 32'h1f5504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1889   :   assert (rdbk == 32'h2460ef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1890   :   assert (rdbk == 32'hf26aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1891   :   assert (rdbk == 32'h429ea1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1892   :   assert (rdbk == 32'h6f39e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1893   :   assert (rdbk == 32'h17a924) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1894   :   assert (rdbk == 32'h590be8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1895   :   assert (rdbk == 32'h6afecd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1896   :   assert (rdbk == 32'h10abcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1897   :   assert (rdbk == 32'hb1493) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1898   :   assert (rdbk == 32'h241345) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1899   :   assert (rdbk == 32'h681684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1900   :   assert (rdbk == 32'h449a89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1901   :   assert (rdbk == 32'h39b474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1902   :   assert (rdbk == 32'h4a93aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1903   :   assert (rdbk == 32'h409e0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1904   :   assert (rdbk == 32'h3924b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1905   :   assert (rdbk == 32'h26ff4d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1906   :   assert (rdbk == 32'h4d07cd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1907   :   assert (rdbk == 32'h60d18f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1908   :   assert (rdbk == 32'h4a837f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1909   :   assert (rdbk == 32'h40d247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1910   :   assert (rdbk == 32'h632c96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1911   :   assert (rdbk == 32'h1acf80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1912   :   assert (rdbk == 32'h7f21bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1913   :   assert (rdbk == 32'h20237b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1914   :   assert (rdbk == 32'h5ba0e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1915   :   assert (rdbk == 32'h37e0dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1916   :   assert (rdbk == 32'h5cae31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1917   :   assert (rdbk == 32'h1b17b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1918   :   assert (rdbk == 32'h1deef9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1919   :   assert (rdbk == 32'h495e78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1920   :   assert (rdbk == 32'h331621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1921   :   assert (rdbk == 32'h1bb646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1922   :   assert (rdbk == 32'h38bd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1923   :   assert (rdbk == 32'h30a029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1924   :   assert (rdbk == 32'hc9eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1925   :   assert (rdbk == 32'haab7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1926   :   assert (rdbk == 32'h193e8c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1927   :   assert (rdbk == 32'h4096fe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1928   :   assert (rdbk == 32'h3ad5ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1929   :   assert (rdbk == 32'h252618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1930   :   assert (rdbk == 32'h36969d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1931   :   assert (rdbk == 32'h583509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1932   :   assert (rdbk == 32'h74d455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1933   :   assert (rdbk == 32'h4e8062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1934   :   assert (rdbk == 32'h4c121b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1935   :   assert (rdbk == 32'h45b9eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1936   :   assert (rdbk == 32'h66311f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1937   :   assert (rdbk == 32'hb1d7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1938   :   assert (rdbk == 32'h536a05) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1939   :   assert (rdbk == 32'h39f270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1940   :   assert (rdbk == 32'hf7e74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1941   :   assert (rdbk == 32'h535102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1942   :   assert (rdbk == 32'h16ae1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1943   :   assert (rdbk == 32'h59a4fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1944   :   assert (rdbk == 32'h47536a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1945   :   assert (rdbk == 32'h25dfe9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1946   :   assert (rdbk == 32'h7724ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1947   :   assert (rdbk == 32'h612c25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1948   :   assert (rdbk == 32'h6ecf13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1949   :   assert (rdbk == 32'h15d960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1950   :   assert (rdbk == 32'h2b7338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1951   :   assert (rdbk == 32'h70f401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1952   :   assert (rdbk == 32'h4cc983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1953   :   assert (rdbk == 32'h98082) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1954   :   assert (rdbk == 32'h2abb7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1955   :   assert (rdbk == 32'h1c3be8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1956   :   assert (rdbk == 32'h3a1ab4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1957   :   assert (rdbk == 32'h6c5a33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1958   :   assert (rdbk == 32'h11e0f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1959   :   assert (rdbk == 32'h5522f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1960   :   assert (rdbk == 32'h6171b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1961   :   assert (rdbk == 32'h23e943) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1962   :   assert (rdbk == 32'h720537) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1963   :   assert (rdbk == 32'h606bb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1964   :   assert (rdbk == 32'he4f98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1965   :   assert (rdbk == 32'h1a6fbb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1966   :   assert (rdbk == 32'h62f4f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1967   :   assert (rdbk == 32'h25dcfe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1968   :   assert (rdbk == 32'h572fff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1969   :   assert (rdbk == 32'h3e42c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1970   :   assert (rdbk == 32'h206b76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1971   :   assert (rdbk == 32'h6fb513) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1972   :   assert (rdbk == 32'h413ff1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1973   :   assert (rdbk == 32'h61141c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1974   :   assert (rdbk == 32'h4112cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1975   :   assert (rdbk == 32'h133028) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1976   :   assert (rdbk == 32'h50da4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1977   :   assert (rdbk == 32'h689df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1978   :   assert (rdbk == 32'h7802fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1979   :   assert (rdbk == 32'hce661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1980   :   assert (rdbk == 32'h4deccc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1981   :   assert (rdbk == 32'h547fd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1982   :   assert (rdbk == 32'h741641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1983   :   assert (rdbk == 32'h372421) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1984   :   assert (rdbk == 32'h793961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1985   :   assert (rdbk == 32'h61c627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1986   :   assert (rdbk == 32'h115bb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1987   :   assert (rdbk == 32'h69e031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1988   :   assert (rdbk == 32'h2adc3e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1989   :   assert (rdbk == 32'h7797ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1990   :   assert (rdbk == 32'h29f8a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1991   :   assert (rdbk == 32'h33ffe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1992   :   assert (rdbk == 32'h66d4b2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1993   :   assert (rdbk == 32'h6a4c59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1994   :   assert (rdbk == 32'h71524d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1995   :   assert (rdbk == 32'h5e2566) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1996   :   assert (rdbk == 32'h34ff32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1997   :   assert (rdbk == 32'h761811) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1998   :   assert (rdbk == 32'h143d40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	1999   :   assert (rdbk == 32'hcca8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2000   :   assert (rdbk == 32'h7487f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2001   :   assert (rdbk == 32'h6c2f97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2002   :   assert (rdbk == 32'h603f48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2003   :   assert (rdbk == 32'h7aa137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2004   :   assert (rdbk == 32'h3d9fb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2005   :   assert (rdbk == 32'h28f84e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2006   :   assert (rdbk == 32'h6fe0b1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2007   :   assert (rdbk == 32'h42e32c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2008   :   assert (rdbk == 32'h141b6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2009   :   assert (rdbk == 32'h4b08ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2010   :   assert (rdbk == 32'h53b6db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2011   :   assert (rdbk == 32'h76cfbb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2012   :   assert (rdbk == 32'hd7a02) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2013   :   assert (rdbk == 32'h219cac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2014   :   assert (rdbk == 32'h1c8e0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2015   :   assert (rdbk == 32'h53914e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2016   :   assert (rdbk == 32'h698dfb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2017   :   assert (rdbk == 32'h3b6a1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2018   :   assert (rdbk == 32'h2f20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2019   :   assert (rdbk == 32'h2e2e22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2020   :   assert (rdbk == 32'h659706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2021   :   assert (rdbk == 32'h1c542c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2022   :   assert (rdbk == 32'h4d4a69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2023   :   assert (rdbk == 32'h219ff5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2024   :   assert (rdbk == 32'h239c75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2025   :   assert (rdbk == 32'h75ffac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2026   :   assert (rdbk == 32'hc53c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2027   :   assert (rdbk == 32'h1a18a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2028   :   assert (rdbk == 32'h183864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2029   :   assert (rdbk == 32'h279ba7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2030   :   assert (rdbk == 32'h632504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2031   :   assert (rdbk == 32'h5aff4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2032   :   assert (rdbk == 32'h5545e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2033   :   assert (rdbk == 32'hf3adb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2034   :   assert (rdbk == 32'h32f6a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2035   :   assert (rdbk == 32'h3ab2b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2036   :   assert (rdbk == 32'h79ff31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2037   :   assert (rdbk == 32'h224a7a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2038   :   assert (rdbk == 32'h2e8a4d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2039   :   assert (rdbk == 32'h669681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2040   :   assert (rdbk == 32'h515a6b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2041   :   assert (rdbk == 32'h72f9a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2042   :   assert (rdbk == 32'h67a187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2043   :   assert (rdbk == 32'h156d58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2044   :   assert (rdbk == 32'h6f1842) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2045   :   assert (rdbk == 32'h595df1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2046   :   assert (rdbk == 32'h16f577) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2047   :   assert (rdbk == 32'h2108eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h200
	2048   :   assert (rdbk == 32'h40489d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2049   :   assert (rdbk == 32'h56706a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2050   :   assert (rdbk == 32'h6c155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2051   :   assert (rdbk == 32'h7e3f60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2052   :   assert (rdbk == 32'h6bdf21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2053   :   assert (rdbk == 32'h3426f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2054   :   assert (rdbk == 32'h5d3f2e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2055   :   assert (rdbk == 32'h79ac73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2056   :   assert (rdbk == 32'h72d330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2057   :   assert (rdbk == 32'h7b045f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2058   :   assert (rdbk == 32'h53f5b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2059   :   assert (rdbk == 32'h168299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2060   :   assert (rdbk == 32'h7c1633) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2061   :   assert (rdbk == 32'h50577d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2062   :   assert (rdbk == 32'h9cf99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2063   :   assert (rdbk == 32'h2b3fa1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2064   :   assert (rdbk == 32'h22f060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2065   :   assert (rdbk == 32'h133256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2066   :   assert (rdbk == 32'h22e473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2067   :   assert (rdbk == 32'h372fb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2068   :   assert (rdbk == 32'h435e56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2069   :   assert (rdbk == 32'h5ba253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2070   :   assert (rdbk == 32'h6355e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2071   :   assert (rdbk == 32'h2a0a97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2072   :   assert (rdbk == 32'h2166cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2073   :   assert (rdbk == 32'h20424c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2074   :   assert (rdbk == 32'h4d2ffd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2075   :   assert (rdbk == 32'h1ee716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2076   :   assert (rdbk == 32'h76b4f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2077   :   assert (rdbk == 32'h172c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2078   :   assert (rdbk == 32'h354a2f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2079   :   assert (rdbk == 32'h2b4ac4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2080   :   assert (rdbk == 32'h7e7926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2081   :   assert (rdbk == 32'h954d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2082   :   assert (rdbk == 32'h6dccf2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2083   :   assert (rdbk == 32'had817) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2084   :   assert (rdbk == 32'h539cf1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2085   :   assert (rdbk == 32'h297d00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2086   :   assert (rdbk == 32'h706391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2087   :   assert (rdbk == 32'h53172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2088   :   assert (rdbk == 32'h2f1570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2089   :   assert (rdbk == 32'h4f0293) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2090   :   assert (rdbk == 32'h31a567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2091   :   assert (rdbk == 32'h56099e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2092   :   assert (rdbk == 32'h59998a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2093   :   assert (rdbk == 32'h51620e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2094   :   assert (rdbk == 32'h561523) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2095   :   assert (rdbk == 32'h1badad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2096   :   assert (rdbk == 32'h4ccf16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2097   :   assert (rdbk == 32'h46b045) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2098   :   assert (rdbk == 32'ha2a3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2099   :   assert (rdbk == 32'h560583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2100   :   assert (rdbk == 32'h4f79af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2101   :   assert (rdbk == 32'h743c23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2102   :   assert (rdbk == 32'h43cc4f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2103   :   assert (rdbk == 32'h700230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2104   :   assert (rdbk == 32'h6f4836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2105   :   assert (rdbk == 32'h28a991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2106   :   assert (rdbk == 32'h3bb664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2107   :   assert (rdbk == 32'h3fef3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2108   :   assert (rdbk == 32'h2abad7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2109   :   assert (rdbk == 32'h9f9ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2110   :   assert (rdbk == 32'h698b5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2111   :   assert (rdbk == 32'h410766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2112   :   assert (rdbk == 32'h30b1e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2113   :   assert (rdbk == 32'h15d87b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2114   :   assert (rdbk == 32'h14d2d9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2115   :   assert (rdbk == 32'h6d8da2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2116   :   assert (rdbk == 32'h476446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2117   :   assert (rdbk == 32'h7bf5b2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2118   :   assert (rdbk == 32'h70f875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2119   :   assert (rdbk == 32'h792cce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2120   :   assert (rdbk == 32'h23a50e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2121   :   assert (rdbk == 32'hbf374) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2122   :   assert (rdbk == 32'h3ffc6a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2123   :   assert (rdbk == 32'h30646a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2124   :   assert (rdbk == 32'h1b154e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2125   :   assert (rdbk == 32'h6325fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2126   :   assert (rdbk == 32'h137e62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2127   :   assert (rdbk == 32'h7dc057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2128   :   assert (rdbk == 32'h1739dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2129   :   assert (rdbk == 32'h6a2422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2130   :   assert (rdbk == 32'h113c55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2131   :   assert (rdbk == 32'h6a0098) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2132   :   assert (rdbk == 32'h4aa52c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2133   :   assert (rdbk == 32'h5cec6b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2134   :   assert (rdbk == 32'h70b138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2135   :   assert (rdbk == 32'h2810d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2136   :   assert (rdbk == 32'h179e3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2137   :   assert (rdbk == 32'h265f7b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2138   :   assert (rdbk == 32'h352561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2139   :   assert (rdbk == 32'h291e5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2140   :   assert (rdbk == 32'h5fb740) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2141   :   assert (rdbk == 32'h202c9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2142   :   assert (rdbk == 32'hbea1a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2143   :   assert (rdbk == 32'h2f7add) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2144   :   assert (rdbk == 32'h6a6bb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2145   :   assert (rdbk == 32'h1161d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2146   :   assert (rdbk == 32'h2754cd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2147   :   assert (rdbk == 32'h50157e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2148   :   assert (rdbk == 32'h6f3934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2149   :   assert (rdbk == 32'h31abd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2150   :   assert (rdbk == 32'h6fad67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2151   :   assert (rdbk == 32'h2ee5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2152   :   assert (rdbk == 32'h52b28e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2153   :   assert (rdbk == 32'h45881e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2154   :   assert (rdbk == 32'h428fbd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2155   :   assert (rdbk == 32'h1a75a4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2156   :   assert (rdbk == 32'h3fb8d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2157   :   assert (rdbk == 32'h349f3e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2158   :   assert (rdbk == 32'h2f8b0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2159   :   assert (rdbk == 32'h717254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2160   :   assert (rdbk == 32'h694b3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2161   :   assert (rdbk == 32'h701380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2162   :   assert (rdbk == 32'h24fc5e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2163   :   assert (rdbk == 32'h3909ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2164   :   assert (rdbk == 32'h2d27bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2165   :   assert (rdbk == 32'h265e07) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2166   :   assert (rdbk == 32'h57ea68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2167   :   assert (rdbk == 32'h408b93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2168   :   assert (rdbk == 32'h3388a1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2169   :   assert (rdbk == 32'h67dfbb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2170   :   assert (rdbk == 32'h37e9b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2171   :   assert (rdbk == 32'h17f13f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2172   :   assert (rdbk == 32'h36dc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2173   :   assert (rdbk == 32'h52050f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2174   :   assert (rdbk == 32'h289f6d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2175   :   assert (rdbk == 32'hbf156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2176   :   assert (rdbk == 32'h49c26b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2177   :   assert (rdbk == 32'h133956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2178   :   assert (rdbk == 32'h655d7a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2179   :   assert (rdbk == 32'h677b1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2180   :   assert (rdbk == 32'h24afd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2181   :   assert (rdbk == 32'h53d930) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2182   :   assert (rdbk == 32'h1248a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2183   :   assert (rdbk == 32'h3186df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2184   :   assert (rdbk == 32'h233960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2185   :   assert (rdbk == 32'h5d6d6c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2186   :   assert (rdbk == 32'h2b0750) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2187   :   assert (rdbk == 32'h331bde) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2188   :   assert (rdbk == 32'h5c5c39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2189   :   assert (rdbk == 32'h4064ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2190   :   assert (rdbk == 32'h6bf006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2191   :   assert (rdbk == 32'h7de384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2192   :   assert (rdbk == 32'h2a0aef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2193   :   assert (rdbk == 32'h6ab163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2194   :   assert (rdbk == 32'h12ba0e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2195   :   assert (rdbk == 32'h14677f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2196   :   assert (rdbk == 32'h3f1e89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2197   :   assert (rdbk == 32'h1a842e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2198   :   assert (rdbk == 32'h42d7e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2199   :   assert (rdbk == 32'h685011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2200   :   assert (rdbk == 32'h66e287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2201   :   assert (rdbk == 32'hab36a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2202   :   assert (rdbk == 32'h372b9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2203   :   assert (rdbk == 32'h75d81a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2204   :   assert (rdbk == 32'h499b90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2205   :   assert (rdbk == 32'h5b60cd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2206   :   assert (rdbk == 32'h4fa62a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2207   :   assert (rdbk == 32'h5344e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2208   :   assert (rdbk == 32'h6b643f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2209   :   assert (rdbk == 32'h4aa717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2210   :   assert (rdbk == 32'h42f5a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2211   :   assert (rdbk == 32'h1187e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2212   :   assert (rdbk == 32'h41ed7c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2213   :   assert (rdbk == 32'h68bc44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2214   :   assert (rdbk == 32'h10bf0a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2215   :   assert (rdbk == 32'h71f2a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2216   :   assert (rdbk == 32'h126eeb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2217   :   assert (rdbk == 32'hc2b45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2218   :   assert (rdbk == 32'h1ec453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2219   :   assert (rdbk == 32'hf26cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2220   :   assert (rdbk == 32'h688045) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2221   :   assert (rdbk == 32'h1f4428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2222   :   assert (rdbk == 32'h42cadf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2223   :   assert (rdbk == 32'h7fb350) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2224   :   assert (rdbk == 32'h6da886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2225   :   assert (rdbk == 32'h610405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2226   :   assert (rdbk == 32'h7c0ff1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2227   :   assert (rdbk == 32'h3af4d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2228   :   assert (rdbk == 32'h6f2e00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2229   :   assert (rdbk == 32'h2a48d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2230   :   assert (rdbk == 32'h213ad0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2231   :   assert (rdbk == 32'h1d84b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2232   :   assert (rdbk == 32'h3dd3dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2233   :   assert (rdbk == 32'h4d3392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2234   :   assert (rdbk == 32'h3f0cb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2235   :   assert (rdbk == 32'h45d9e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2236   :   assert (rdbk == 32'h370fe8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2237   :   assert (rdbk == 32'h1ac68c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2238   :   assert (rdbk == 32'h1923bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2239   :   assert (rdbk == 32'h59f72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2240   :   assert (rdbk == 32'h6caaa2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2241   :   assert (rdbk == 32'h4f0a0c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2242   :   assert (rdbk == 32'h7da6a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2243   :   assert (rdbk == 32'hc2753) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2244   :   assert (rdbk == 32'h6fd4d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2245   :   assert (rdbk == 32'h7ac4d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2246   :   assert (rdbk == 32'h17dffe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2247   :   assert (rdbk == 32'h3efce8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2248   :   assert (rdbk == 32'h209d47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2249   :   assert (rdbk == 32'h609896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2250   :   assert (rdbk == 32'h62e126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2251   :   assert (rdbk == 32'h7a639a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2252   :   assert (rdbk == 32'hbc22b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2253   :   assert (rdbk == 32'h68803b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2254   :   assert (rdbk == 32'h22ac2a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2255   :   assert (rdbk == 32'h11ab31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2256   :   assert (rdbk == 32'h6bbc37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2257   :   assert (rdbk == 32'h4a5dcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2258   :   assert (rdbk == 32'h73f077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2259   :   assert (rdbk == 32'h6cfbf1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2260   :   assert (rdbk == 32'h3e60c6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2261   :   assert (rdbk == 32'h510911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2262   :   assert (rdbk == 32'h73fa99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2263   :   assert (rdbk == 32'h27a783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2264   :   assert (rdbk == 32'h6bb6b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2265   :   assert (rdbk == 32'h57077e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2266   :   assert (rdbk == 32'h50305e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2267   :   assert (rdbk == 32'h570d1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2268   :   assert (rdbk == 32'h7a465a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2269   :   assert (rdbk == 32'h403742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2270   :   assert (rdbk == 32'h58fec7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2271   :   assert (rdbk == 32'h70d39a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2272   :   assert (rdbk == 32'h4ca1ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2273   :   assert (rdbk == 32'h288302) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2274   :   assert (rdbk == 32'h16bdd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2275   :   assert (rdbk == 32'h57ec41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2276   :   assert (rdbk == 32'h2edeb1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2277   :   assert (rdbk == 32'h3b90ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2278   :   assert (rdbk == 32'h175d4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2279   :   assert (rdbk == 32'h35137f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2280   :   assert (rdbk == 32'h562616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2281   :   assert (rdbk == 32'h5330b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2282   :   assert (rdbk == 32'h1a3383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2283   :   assert (rdbk == 32'h43d1d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2284   :   assert (rdbk == 32'h7a22c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2285   :   assert (rdbk == 32'h29c3cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2286   :   assert (rdbk == 32'h277d1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2287   :   assert (rdbk == 32'h524e4e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2288   :   assert (rdbk == 32'hd70b1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2289   :   assert (rdbk == 32'h1b7eb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2290   :   assert (rdbk == 32'h4a7fd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2291   :   assert (rdbk == 32'h47d773) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2292   :   assert (rdbk == 32'h7b0f73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2293   :   assert (rdbk == 32'h53597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2294   :   assert (rdbk == 32'h74475f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2295   :   assert (rdbk == 32'h1ff71b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2296   :   assert (rdbk == 32'h70df20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2297   :   assert (rdbk == 32'h68dbd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2298   :   assert (rdbk == 32'h210d52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2299   :   assert (rdbk == 32'h1bfa0a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2300   :   assert (rdbk == 32'h7d97c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2301   :   assert (rdbk == 32'h145e6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2302   :   assert (rdbk == 32'h705441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2303   :   assert (rdbk == 32'h3c01cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h201
	2304   :   assert (rdbk == 32'h4de661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2305   :   assert (rdbk == 32'h3bbae6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2306   :   assert (rdbk == 32'h45f5d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2307   :   assert (rdbk == 32'h513a65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2308   :   assert (rdbk == 32'h5bcfd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2309   :   assert (rdbk == 32'ha1636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2310   :   assert (rdbk == 32'h664b98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2311   :   assert (rdbk == 32'h44c09) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2312   :   assert (rdbk == 32'h451266) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2313   :   assert (rdbk == 32'h6d7dea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2314   :   assert (rdbk == 32'h65abaf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2315   :   assert (rdbk == 32'h327702) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2316   :   assert (rdbk == 32'hb0160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2317   :   assert (rdbk == 32'h3b7254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2318   :   assert (rdbk == 32'h3655dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2319   :   assert (rdbk == 32'h3d58d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2320   :   assert (rdbk == 32'h63067a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2321   :   assert (rdbk == 32'h12f5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2322   :   assert (rdbk == 32'h2680c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2323   :   assert (rdbk == 32'h7cbaeb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2324   :   assert (rdbk == 32'h579263) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2325   :   assert (rdbk == 32'h1626d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2326   :   assert (rdbk == 32'hf7251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2327   :   assert (rdbk == 32'h23629) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2328   :   assert (rdbk == 32'habb54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2329   :   assert (rdbk == 32'h16272a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2330   :   assert (rdbk == 32'h157218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2331   :   assert (rdbk == 32'hac46f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2332   :   assert (rdbk == 32'h6acb5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2333   :   assert (rdbk == 32'h7b359f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2334   :   assert (rdbk == 32'h6c7626) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2335   :   assert (rdbk == 32'h201aaf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2336   :   assert (rdbk == 32'h5451e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2337   :   assert (rdbk == 32'h399084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2338   :   assert (rdbk == 32'h7694ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2339   :   assert (rdbk == 32'h43efc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2340   :   assert (rdbk == 32'h7ba88c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2341   :   assert (rdbk == 32'h269688) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2342   :   assert (rdbk == 32'h739427) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2343   :   assert (rdbk == 32'h7bd59b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2344   :   assert (rdbk == 32'h38ceac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2345   :   assert (rdbk == 32'h6497e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2346   :   assert (rdbk == 32'h435a67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2347   :   assert (rdbk == 32'h3ccc0c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2348   :   assert (rdbk == 32'h10d3ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2349   :   assert (rdbk == 32'h1d0691) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2350   :   assert (rdbk == 32'h3040e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2351   :   assert (rdbk == 32'h5ceef3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2352   :   assert (rdbk == 32'h35e99a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2353   :   assert (rdbk == 32'h5af390) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2354   :   assert (rdbk == 32'h399e17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2355   :   assert (rdbk == 32'h2d3f4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2356   :   assert (rdbk == 32'h6f4aa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2357   :   assert (rdbk == 32'h45a528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2358   :   assert (rdbk == 32'h4fc65b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2359   :   assert (rdbk == 32'h37313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2360   :   assert (rdbk == 32'h3b9dd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2361   :   assert (rdbk == 32'h24efe9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2362   :   assert (rdbk == 32'h2e22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2363   :   assert (rdbk == 32'h76605c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2364   :   assert (rdbk == 32'h7d5ef6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2365   :   assert (rdbk == 32'h77a0bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2366   :   assert (rdbk == 32'h27c211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2367   :   assert (rdbk == 32'h3d7dc4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2368   :   assert (rdbk == 32'h216b02) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2369   :   assert (rdbk == 32'h1d5c83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2370   :   assert (rdbk == 32'h660ebf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2371   :   assert (rdbk == 32'h484252) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2372   :   assert (rdbk == 32'h46230d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2373   :   assert (rdbk == 32'h3549df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2374   :   assert (rdbk == 32'h7da53c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2375   :   assert (rdbk == 32'h545490) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2376   :   assert (rdbk == 32'h230243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2377   :   assert (rdbk == 32'hb1ffe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2378   :   assert (rdbk == 32'h1ea9f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2379   :   assert (rdbk == 32'hf9271) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2380   :   assert (rdbk == 32'h38fff7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2381   :   assert (rdbk == 32'h43442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2382   :   assert (rdbk == 32'h73cc93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2383   :   assert (rdbk == 32'h557ec2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2384   :   assert (rdbk == 32'h69f2a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2385   :   assert (rdbk == 32'h5739e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2386   :   assert (rdbk == 32'hafccb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2387   :   assert (rdbk == 32'h26b172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2388   :   assert (rdbk == 32'h51dd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2389   :   assert (rdbk == 32'h55b72a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2390   :   assert (rdbk == 32'h5b1550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2391   :   assert (rdbk == 32'h796bed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2392   :   assert (rdbk == 32'h186eb8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2393   :   assert (rdbk == 32'h2737c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2394   :   assert (rdbk == 32'h72b8d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2395   :   assert (rdbk == 32'h270dab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2396   :   assert (rdbk == 32'h691d14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2397   :   assert (rdbk == 32'h442c89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2398   :   assert (rdbk == 32'h18a6d9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2399   :   assert (rdbk == 32'h60e193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2400   :   assert (rdbk == 32'h2b4623) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2401   :   assert (rdbk == 32'h583825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2402   :   assert (rdbk == 32'h177551) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2403   :   assert (rdbk == 32'h2b091c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2404   :   assert (rdbk == 32'h3cfce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2405   :   assert (rdbk == 32'h7ec899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2406   :   assert (rdbk == 32'h4c8498) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2407   :   assert (rdbk == 32'h14a804) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2408   :   assert (rdbk == 32'h27fb70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2409   :   assert (rdbk == 32'h6aae5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2410   :   assert (rdbk == 32'h6b28a1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2411   :   assert (rdbk == 32'h6f5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2412   :   assert (rdbk == 32'h16a9ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2413   :   assert (rdbk == 32'h5b0e30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2414   :   assert (rdbk == 32'h7428e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2415   :   assert (rdbk == 32'h10534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2416   :   assert (rdbk == 32'h7b78cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2417   :   assert (rdbk == 32'h76c933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2418   :   assert (rdbk == 32'h51cf01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2419   :   assert (rdbk == 32'h2726a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2420   :   assert (rdbk == 32'h11be01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2421   :   assert (rdbk == 32'h79b80c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2422   :   assert (rdbk == 32'h5e34d9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2423   :   assert (rdbk == 32'h3141f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2424   :   assert (rdbk == 32'h161378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2425   :   assert (rdbk == 32'h116aa7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2426   :   assert (rdbk == 32'h64543a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2427   :   assert (rdbk == 32'h13fc26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2428   :   assert (rdbk == 32'h79c3f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2429   :   assert (rdbk == 32'h28b947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2430   :   assert (rdbk == 32'h73bed0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2431   :   assert (rdbk == 32'h628f1f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2432   :   assert (rdbk == 32'h6fde2b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2433   :   assert (rdbk == 32'h5a68e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2434   :   assert (rdbk == 32'h1a0f36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2435   :   assert (rdbk == 32'h689cea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2436   :   assert (rdbk == 32'h5e0fc7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2437   :   assert (rdbk == 32'h4a4222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2438   :   assert (rdbk == 32'h513a49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2439   :   assert (rdbk == 32'h773d5e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2440   :   assert (rdbk == 32'h41f052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2441   :   assert (rdbk == 32'h348e30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2442   :   assert (rdbk == 32'h34d000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2443   :   assert (rdbk == 32'h50293f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2444   :   assert (rdbk == 32'h6703f4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2445   :   assert (rdbk == 32'h55fa64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2446   :   assert (rdbk == 32'h477d0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2447   :   assert (rdbk == 32'h3d78fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2448   :   assert (rdbk == 32'h4191fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2449   :   assert (rdbk == 32'h34fe07) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2450   :   assert (rdbk == 32'h6f382d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2451   :   assert (rdbk == 32'hf9e82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2452   :   assert (rdbk == 32'h306bfb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2453   :   assert (rdbk == 32'h3f4a9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2454   :   assert (rdbk == 32'h47a33a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2455   :   assert (rdbk == 32'h1afa6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2456   :   assert (rdbk == 32'h2be5ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2457   :   assert (rdbk == 32'h4de42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2458   :   assert (rdbk == 32'h7c7d1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2459   :   assert (rdbk == 32'h6f0ae1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2460   :   assert (rdbk == 32'h688f9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2461   :   assert (rdbk == 32'h80a7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2462   :   assert (rdbk == 32'h4154e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2463   :   assert (rdbk == 32'h272303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2464   :   assert (rdbk == 32'h29e35c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2465   :   assert (rdbk == 32'h5ea838) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2466   :   assert (rdbk == 32'h1a29d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2467   :   assert (rdbk == 32'h5dc204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2468   :   assert (rdbk == 32'h451978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2469   :   assert (rdbk == 32'h25340b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2470   :   assert (rdbk == 32'hced2d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2471   :   assert (rdbk == 32'h59d5c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2472   :   assert (rdbk == 32'h8d287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2473   :   assert (rdbk == 32'h58e5c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2474   :   assert (rdbk == 32'h6dc5d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2475   :   assert (rdbk == 32'h6ea0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2476   :   assert (rdbk == 32'h1d0a60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2477   :   assert (rdbk == 32'h6e4504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2478   :   assert (rdbk == 32'h51d43b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2479   :   assert (rdbk == 32'h55b7cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2480   :   assert (rdbk == 32'h2bc3a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2481   :   assert (rdbk == 32'h2c81d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2482   :   assert (rdbk == 32'h4e0beb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2483   :   assert (rdbk == 32'h4c00df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2484   :   assert (rdbk == 32'h495763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2485   :   assert (rdbk == 32'h6ac141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2486   :   assert (rdbk == 32'h414f66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2487   :   assert (rdbk == 32'h582783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2488   :   assert (rdbk == 32'h71123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2489   :   assert (rdbk == 32'h733ff3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2490   :   assert (rdbk == 32'h7cc757) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2491   :   assert (rdbk == 32'h671322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2492   :   assert (rdbk == 32'hd09) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2493   :   assert (rdbk == 32'h65ebb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2494   :   assert (rdbk == 32'h72ce92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2495   :   assert (rdbk == 32'h30b55f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2496   :   assert (rdbk == 32'h7f086c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2497   :   assert (rdbk == 32'h645461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2498   :   assert (rdbk == 32'h60219d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2499   :   assert (rdbk == 32'h7c3c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2500   :   assert (rdbk == 32'h2ef789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2501   :   assert (rdbk == 32'h584278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2502   :   assert (rdbk == 32'h158b0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2503   :   assert (rdbk == 32'h158518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2504   :   assert (rdbk == 32'h6d12c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2505   :   assert (rdbk == 32'h16f21d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2506   :   assert (rdbk == 32'h6a5af6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2507   :   assert (rdbk == 32'h325c30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2508   :   assert (rdbk == 32'h19da67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2509   :   assert (rdbk == 32'h54abe2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2510   :   assert (rdbk == 32'h695b9c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2511   :   assert (rdbk == 32'h3c9b1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2512   :   assert (rdbk == 32'h244057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2513   :   assert (rdbk == 32'h7019cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2514   :   assert (rdbk == 32'h4a82d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2515   :   assert (rdbk == 32'h601469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2516   :   assert (rdbk == 32'h7c418f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2517   :   assert (rdbk == 32'h3daddd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2518   :   assert (rdbk == 32'h245cfb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2519   :   assert (rdbk == 32'h75f571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2520   :   assert (rdbk == 32'h77092a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2521   :   assert (rdbk == 32'h3e2a4b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2522   :   assert (rdbk == 32'h57d2a4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2523   :   assert (rdbk == 32'h525e49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2524   :   assert (rdbk == 32'h5562a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2525   :   assert (rdbk == 32'h448d9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2526   :   assert (rdbk == 32'h60522e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2527   :   assert (rdbk == 32'h1d2efb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2528   :   assert (rdbk == 32'h5967ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2529   :   assert (rdbk == 32'h4791e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2530   :   assert (rdbk == 32'h7e5f3a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2531   :   assert (rdbk == 32'h5dc1a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2532   :   assert (rdbk == 32'h7c9f49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2533   :   assert (rdbk == 32'h2b84fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2534   :   assert (rdbk == 32'h27c06d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2535   :   assert (rdbk == 32'h7fd425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2536   :   assert (rdbk == 32'h2bec5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2537   :   assert (rdbk == 32'h7281c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2538   :   assert (rdbk == 32'h1f6659) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2539   :   assert (rdbk == 32'h2c12c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2540   :   assert (rdbk == 32'h8f3d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2541   :   assert (rdbk == 32'h177833) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2542   :   assert (rdbk == 32'h200339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2543   :   assert (rdbk == 32'h1325d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2544   :   assert (rdbk == 32'h1b911a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2545   :   assert (rdbk == 32'hab67b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2546   :   assert (rdbk == 32'h7e6ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2547   :   assert (rdbk == 32'h71859c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2548   :   assert (rdbk == 32'h68bd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2549   :   assert (rdbk == 32'h5cef94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2550   :   assert (rdbk == 32'h710732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2551   :   assert (rdbk == 32'hdff96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2552   :   assert (rdbk == 32'h1b0bf2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2553   :   assert (rdbk == 32'h4e0109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2554   :   assert (rdbk == 32'h7784be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2555   :   assert (rdbk == 32'h3426a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2556   :   assert (rdbk == 32'h1c68b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2557   :   assert (rdbk == 32'h3d75f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2558   :   assert (rdbk == 32'h2cd9c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2559   :   assert (rdbk == 32'h1c5c72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h202
	2560   :   assert (rdbk == 32'h46f21d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2561   :   assert (rdbk == 32'h7fcdc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2562   :   assert (rdbk == 32'h44f946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2563   :   assert (rdbk == 32'h51fee6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2564   :   assert (rdbk == 32'h6bf167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2565   :   assert (rdbk == 32'hcb3eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2566   :   assert (rdbk == 32'h51338a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2567   :   assert (rdbk == 32'h6aecc2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2568   :   assert (rdbk == 32'h38295f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2569   :   assert (rdbk == 32'h13e657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2570   :   assert (rdbk == 32'h54e3d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2571   :   assert (rdbk == 32'h3487bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2572   :   assert (rdbk == 32'h32f2f9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2573   :   assert (rdbk == 32'h1c2df6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2574   :   assert (rdbk == 32'h6ab2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2575   :   assert (rdbk == 32'h586e3b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2576   :   assert (rdbk == 32'h297e8d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2577   :   assert (rdbk == 32'h18a390) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2578   :   assert (rdbk == 32'h36ea96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2579   :   assert (rdbk == 32'hecbd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2580   :   assert (rdbk == 32'h6efe93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2581   :   assert (rdbk == 32'h5932d9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2582   :   assert (rdbk == 32'h66a318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2583   :   assert (rdbk == 32'h1b8057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2584   :   assert (rdbk == 32'h5aba48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2585   :   assert (rdbk == 32'h3de81d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2586   :   assert (rdbk == 32'h14413c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2587   :   assert (rdbk == 32'h184c43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2588   :   assert (rdbk == 32'h39cd92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2589   :   assert (rdbk == 32'h6ca825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2590   :   assert (rdbk == 32'h1c382f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2591   :   assert (rdbk == 32'h28ac63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2592   :   assert (rdbk == 32'ha9fb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2593   :   assert (rdbk == 32'h2f353d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2594   :   assert (rdbk == 32'h76fb60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2595   :   assert (rdbk == 32'h7dcf61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2596   :   assert (rdbk == 32'h6b426c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2597   :   assert (rdbk == 32'h3974e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2598   :   assert (rdbk == 32'h76d213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2599   :   assert (rdbk == 32'h596a19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2600   :   assert (rdbk == 32'h624ea7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2601   :   assert (rdbk == 32'h7258b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2602   :   assert (rdbk == 32'h75d8ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2603   :   assert (rdbk == 32'h28ca69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2604   :   assert (rdbk == 32'h7b08df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2605   :   assert (rdbk == 32'h170411) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2606   :   assert (rdbk == 32'h7fecc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2607   :   assert (rdbk == 32'hef694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2608   :   assert (rdbk == 32'h7abdfa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2609   :   assert (rdbk == 32'h4e52d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2610   :   assert (rdbk == 32'h4adb31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2611   :   assert (rdbk == 32'h7cf679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2612   :   assert (rdbk == 32'h285fef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2613   :   assert (rdbk == 32'h56d22e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2614   :   assert (rdbk == 32'h16e21f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2615   :   assert (rdbk == 32'h1b0ce9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2616   :   assert (rdbk == 32'h223703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2617   :   assert (rdbk == 32'h7cdc21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2618   :   assert (rdbk == 32'h58d46c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2619   :   assert (rdbk == 32'h319024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2620   :   assert (rdbk == 32'h29ed15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2621   :   assert (rdbk == 32'h3335ba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2622   :   assert (rdbk == 32'h44353) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2623   :   assert (rdbk == 32'h3d0d24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2624   :   assert (rdbk == 32'h7e450a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2625   :   assert (rdbk == 32'hd308d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2626   :   assert (rdbk == 32'h4d3179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2627   :   assert (rdbk == 32'h635205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2628   :   assert (rdbk == 32'h7ba8ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2629   :   assert (rdbk == 32'h7978ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2630   :   assert (rdbk == 32'h4e7589) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2631   :   assert (rdbk == 32'h36533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2632   :   assert (rdbk == 32'h753be7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2633   :   assert (rdbk == 32'h12dc9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2634   :   assert (rdbk == 32'h798319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2635   :   assert (rdbk == 32'h641eb6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2636   :   assert (rdbk == 32'h6c6cc4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2637   :   assert (rdbk == 32'h9eabd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2638   :   assert (rdbk == 32'h6131f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2639   :   assert (rdbk == 32'hb0d81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2640   :   assert (rdbk == 32'h47089d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2641   :   assert (rdbk == 32'h2d66c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2642   :   assert (rdbk == 32'h32b1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2643   :   assert (rdbk == 32'h1a0a5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2644   :   assert (rdbk == 32'h61355c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2645   :   assert (rdbk == 32'h16a530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2646   :   assert (rdbk == 32'h78a4f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2647   :   assert (rdbk == 32'h3c6cd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2648   :   assert (rdbk == 32'h400796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2649   :   assert (rdbk == 32'h6a4d00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2650   :   assert (rdbk == 32'h4a5d7c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2651   :   assert (rdbk == 32'h32e7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2652   :   assert (rdbk == 32'h6f7662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2653   :   assert (rdbk == 32'h75c0d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2654   :   assert (rdbk == 32'h551239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2655   :   assert (rdbk == 32'h79cc4f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2656   :   assert (rdbk == 32'h4a7975) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2657   :   assert (rdbk == 32'h52281d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2658   :   assert (rdbk == 32'h574879) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2659   :   assert (rdbk == 32'h6a81d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2660   :   assert (rdbk == 32'h48a13c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2661   :   assert (rdbk == 32'h55b07d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2662   :   assert (rdbk == 32'h21abb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2663   :   assert (rdbk == 32'h747513) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2664   :   assert (rdbk == 32'h46d748) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2665   :   assert (rdbk == 32'h6fac22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2666   :   assert (rdbk == 32'h66b1c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2667   :   assert (rdbk == 32'h3c2b09) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2668   :   assert (rdbk == 32'h3d2610) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2669   :   assert (rdbk == 32'h364528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2670   :   assert (rdbk == 32'h1f0e0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2671   :   assert (rdbk == 32'h497bd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2672   :   assert (rdbk == 32'h1a8f9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2673   :   assert (rdbk == 32'h73543) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2674   :   assert (rdbk == 32'h9eaff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2675   :   assert (rdbk == 32'h48af1e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2676   :   assert (rdbk == 32'h2a49f4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2677   :   assert (rdbk == 32'h7d4fdf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2678   :   assert (rdbk == 32'h464215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2679   :   assert (rdbk == 32'h2ca510) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2680   :   assert (rdbk == 32'h3efa25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2681   :   assert (rdbk == 32'h305756) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2682   :   assert (rdbk == 32'h6a365a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2683   :   assert (rdbk == 32'h60e82e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2684   :   assert (rdbk == 32'h410275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2685   :   assert (rdbk == 32'he4c12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2686   :   assert (rdbk == 32'h20269a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2687   :   assert (rdbk == 32'h6db25a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2688   :   assert (rdbk == 32'h441f3e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2689   :   assert (rdbk == 32'h4bfe29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2690   :   assert (rdbk == 32'h17adbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2691   :   assert (rdbk == 32'h472802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2692   :   assert (rdbk == 32'hc2650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2693   :   assert (rdbk == 32'h40e730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2694   :   assert (rdbk == 32'h3dbe5e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2695   :   assert (rdbk == 32'h4fe5f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2696   :   assert (rdbk == 32'h246f02) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2697   :   assert (rdbk == 32'h2c3066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2698   :   assert (rdbk == 32'h49a5f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2699   :   assert (rdbk == 32'h74ad01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2700   :   assert (rdbk == 32'h22befe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2701   :   assert (rdbk == 32'h213304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2702   :   assert (rdbk == 32'h65aa4c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2703   :   assert (rdbk == 32'h61c9a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2704   :   assert (rdbk == 32'he18ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2705   :   assert (rdbk == 32'h6c7062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2706   :   assert (rdbk == 32'h781f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2707   :   assert (rdbk == 32'h8d911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2708   :   assert (rdbk == 32'h79ac1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2709   :   assert (rdbk == 32'h287945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2710   :   assert (rdbk == 32'h173b3c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2711   :   assert (rdbk == 32'h1c9ea3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2712   :   assert (rdbk == 32'h5ee62f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2713   :   assert (rdbk == 32'h229895) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2714   :   assert (rdbk == 32'h29ebe2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2715   :   assert (rdbk == 32'h38be50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2716   :   assert (rdbk == 32'h5f4209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2717   :   assert (rdbk == 32'h1e5c4d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2718   :   assert (rdbk == 32'h32d6b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2719   :   assert (rdbk == 32'h596dd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2720   :   assert (rdbk == 32'h258d23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2721   :   assert (rdbk == 32'h47c4b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2722   :   assert (rdbk == 32'h4531b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2723   :   assert (rdbk == 32'h38b401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2724   :   assert (rdbk == 32'h4370c3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2725   :   assert (rdbk == 32'h770ea5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2726   :   assert (rdbk == 32'haf40b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2727   :   assert (rdbk == 32'h5b7ef2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2728   :   assert (rdbk == 32'h194529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2729   :   assert (rdbk == 32'hedf67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2730   :   assert (rdbk == 32'h34c121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2731   :   assert (rdbk == 32'h3180c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2732   :   assert (rdbk == 32'h68aac6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2733   :   assert (rdbk == 32'h6ca03d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2734   :   assert (rdbk == 32'h54b899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2735   :   assert (rdbk == 32'h9b7bf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2736   :   assert (rdbk == 32'h1d5bee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2737   :   assert (rdbk == 32'h3b4d25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2738   :   assert (rdbk == 32'h64a686) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2739   :   assert (rdbk == 32'h77c25f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2740   :   assert (rdbk == 32'h40e4af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2741   :   assert (rdbk == 32'h497e36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2742   :   assert (rdbk == 32'h205c24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2743   :   assert (rdbk == 32'h69167c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2744   :   assert (rdbk == 32'h62a9b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2745   :   assert (rdbk == 32'h33d68f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2746   :   assert (rdbk == 32'h327e93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2747   :   assert (rdbk == 32'h6dc88c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2748   :   assert (rdbk == 32'h1d238a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2749   :   assert (rdbk == 32'h7b7d2f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2750   :   assert (rdbk == 32'h1f3549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2751   :   assert (rdbk == 32'h6d00d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2752   :   assert (rdbk == 32'h2f7cb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2753   :   assert (rdbk == 32'h5acaad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2754   :   assert (rdbk == 32'h4831d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2755   :   assert (rdbk == 32'h13013d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2756   :   assert (rdbk == 32'h42b7dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2757   :   assert (rdbk == 32'h4e1874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2758   :   assert (rdbk == 32'h4106e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2759   :   assert (rdbk == 32'h60038c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2760   :   assert (rdbk == 32'h606bad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2761   :   assert (rdbk == 32'haf17d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2762   :   assert (rdbk == 32'h2b11e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2763   :   assert (rdbk == 32'h61eda3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2764   :   assert (rdbk == 32'h20fa3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2765   :   assert (rdbk == 32'hdf828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2766   :   assert (rdbk == 32'h462afb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2767   :   assert (rdbk == 32'hbaa47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2768   :   assert (rdbk == 32'h72bcab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2769   :   assert (rdbk == 32'h43e2df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2770   :   assert (rdbk == 32'h48d43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2771   :   assert (rdbk == 32'h7aae6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2772   :   assert (rdbk == 32'h671a6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2773   :   assert (rdbk == 32'h7b095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2774   :   assert (rdbk == 32'h433ef4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2775   :   assert (rdbk == 32'h65b142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2776   :   assert (rdbk == 32'h13497d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2777   :   assert (rdbk == 32'h1315a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2778   :   assert (rdbk == 32'h5a33bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2779   :   assert (rdbk == 32'h22b793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2780   :   assert (rdbk == 32'h28ee1f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2781   :   assert (rdbk == 32'h54b061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2782   :   assert (rdbk == 32'h61609f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2783   :   assert (rdbk == 32'h4eed04) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2784   :   assert (rdbk == 32'h482354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2785   :   assert (rdbk == 32'haf9b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2786   :   assert (rdbk == 32'h424d47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2787   :   assert (rdbk == 32'h7355b2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2788   :   assert (rdbk == 32'h367ce5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2789   :   assert (rdbk == 32'h312905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2790   :   assert (rdbk == 32'h2b841d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2791   :   assert (rdbk == 32'h56fd89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2792   :   assert (rdbk == 32'h5840ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2793   :   assert (rdbk == 32'h13409c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2794   :   assert (rdbk == 32'h12a122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2795   :   assert (rdbk == 32'h7aa324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2796   :   assert (rdbk == 32'h62d28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2797   :   assert (rdbk == 32'h20adf0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2798   :   assert (rdbk == 32'h8e099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2799   :   assert (rdbk == 32'h73a2e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2800   :   assert (rdbk == 32'h30a2dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2801   :   assert (rdbk == 32'h66338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2802   :   assert (rdbk == 32'h761b28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2803   :   assert (rdbk == 32'h193d55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2804   :   assert (rdbk == 32'h6fb762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2805   :   assert (rdbk == 32'h4e981e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2806   :   assert (rdbk == 32'h37f9a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2807   :   assert (rdbk == 32'h59f9d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2808   :   assert (rdbk == 32'ha444c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2809   :   assert (rdbk == 32'h5bca26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2810   :   assert (rdbk == 32'h55cee0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2811   :   assert (rdbk == 32'h2581f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2812   :   assert (rdbk == 32'h41681a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2813   :   assert (rdbk == 32'h1ef869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2814   :   assert (rdbk == 32'h168565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2815   :   assert (rdbk == 32'h6bafc4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h203
	2816   :   assert (rdbk == 32'h5e8b38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2817   :   assert (rdbk == 32'h47089f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2818   :   assert (rdbk == 32'h798fde) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2819   :   assert (rdbk == 32'h2d523) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2820   :   assert (rdbk == 32'h4fa459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2821   :   assert (rdbk == 32'h689fc1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2822   :   assert (rdbk == 32'h206fe0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2823   :   assert (rdbk == 32'h3ba84a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2824   :   assert (rdbk == 32'h2e90e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2825   :   assert (rdbk == 32'h51a09) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2826   :   assert (rdbk == 32'h66e5d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2827   :   assert (rdbk == 32'h39c6eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2828   :   assert (rdbk == 32'h584c88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2829   :   assert (rdbk == 32'h196e35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2830   :   assert (rdbk == 32'h44c6a9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2831   :   assert (rdbk == 32'h561694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2832   :   assert (rdbk == 32'h6d2e30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2833   :   assert (rdbk == 32'h1758d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2834   :   assert (rdbk == 32'h70706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2835   :   assert (rdbk == 32'h4eac15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2836   :   assert (rdbk == 32'h320dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2837   :   assert (rdbk == 32'h605f23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2838   :   assert (rdbk == 32'h73293) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2839   :   assert (rdbk == 32'h6f738) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2840   :   assert (rdbk == 32'h5c923b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2841   :   assert (rdbk == 32'h492ef2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2842   :   assert (rdbk == 32'h2c1757) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2843   :   assert (rdbk == 32'h4527a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2844   :   assert (rdbk == 32'h6beccb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2845   :   assert (rdbk == 32'h7b946b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2846   :   assert (rdbk == 32'h73f5d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2847   :   assert (rdbk == 32'h7fc206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2848   :   assert (rdbk == 32'h5d0f97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2849   :   assert (rdbk == 32'h2bf70b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2850   :   assert (rdbk == 32'h1715a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2851   :   assert (rdbk == 32'h6ed393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2852   :   assert (rdbk == 32'h357d97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2853   :   assert (rdbk == 32'h300369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2854   :   assert (rdbk == 32'h6efdef) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2855   :   assert (rdbk == 32'h442894) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2856   :   assert (rdbk == 32'h2dd080) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2857   :   assert (rdbk == 32'h7a995e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2858   :   assert (rdbk == 32'h446c85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2859   :   assert (rdbk == 32'h63ee9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2860   :   assert (rdbk == 32'h6ce5a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2861   :   assert (rdbk == 32'h68a78c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2862   :   assert (rdbk == 32'h452c5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2863   :   assert (rdbk == 32'h56f98f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2864   :   assert (rdbk == 32'h212b0c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2865   :   assert (rdbk == 32'h192504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2866   :   assert (rdbk == 32'h474283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2867   :   assert (rdbk == 32'h4fa1c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2868   :   assert (rdbk == 32'h780bd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2869   :   assert (rdbk == 32'h487f7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2870   :   assert (rdbk == 32'h5f6799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2871   :   assert (rdbk == 32'h21e94f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2872   :   assert (rdbk == 32'h2f3a97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2873   :   assert (rdbk == 32'h6b7744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2874   :   assert (rdbk == 32'h34c16c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2875   :   assert (rdbk == 32'h232bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2876   :   assert (rdbk == 32'h57e7c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2877   :   assert (rdbk == 32'h41d027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2878   :   assert (rdbk == 32'h303dd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2879   :   assert (rdbk == 32'h686083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2880   :   assert (rdbk == 32'h501f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2881   :   assert (rdbk == 32'h2dd2c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2882   :   assert (rdbk == 32'h1f3dec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2883   :   assert (rdbk == 32'h589cea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2884   :   assert (rdbk == 32'h225fe3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2885   :   assert (rdbk == 32'h8c135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2886   :   assert (rdbk == 32'h7d0b1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2887   :   assert (rdbk == 32'h5f637f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2888   :   assert (rdbk == 32'h3e7979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2889   :   assert (rdbk == 32'h6ab967) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2890   :   assert (rdbk == 32'h704512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2891   :   assert (rdbk == 32'h4ceb40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2892   :   assert (rdbk == 32'h6eface) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2893   :   assert (rdbk == 32'h38043c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2894   :   assert (rdbk == 32'h336705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2895   :   assert (rdbk == 32'h5c3e48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2896   :   assert (rdbk == 32'h5c6013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2897   :   assert (rdbk == 32'h3b9131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2898   :   assert (rdbk == 32'h327bd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2899   :   assert (rdbk == 32'h58dd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2900   :   assert (rdbk == 32'h291ddc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2901   :   assert (rdbk == 32'ha5df2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2902   :   assert (rdbk == 32'h649b47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2903   :   assert (rdbk == 32'h730c94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2904   :   assert (rdbk == 32'h3467ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2905   :   assert (rdbk == 32'h379768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2906   :   assert (rdbk == 32'h4abc69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2907   :   assert (rdbk == 32'h6ca97f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2908   :   assert (rdbk == 32'h65e8af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2909   :   assert (rdbk == 32'h72a74b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2910   :   assert (rdbk == 32'h23a8d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2911   :   assert (rdbk == 32'h5b31f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2912   :   assert (rdbk == 32'h69f4bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2913   :   assert (rdbk == 32'h66d917) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2914   :   assert (rdbk == 32'h647f1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2915   :   assert (rdbk == 32'h670f68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2916   :   assert (rdbk == 32'hf61dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2917   :   assert (rdbk == 32'h10a2fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2918   :   assert (rdbk == 32'h27dee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2919   :   assert (rdbk == 32'h4d7bd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2920   :   assert (rdbk == 32'hbf6cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2921   :   assert (rdbk == 32'h4a0d9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2922   :   assert (rdbk == 32'h2afd3b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2923   :   assert (rdbk == 32'h76ca8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2924   :   assert (rdbk == 32'h1b4968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2925   :   assert (rdbk == 32'h32195a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2926   :   assert (rdbk == 32'h38bce9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2927   :   assert (rdbk == 32'h740a85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2928   :   assert (rdbk == 32'h16ecda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2929   :   assert (rdbk == 32'h6842fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2930   :   assert (rdbk == 32'h5bf1dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2931   :   assert (rdbk == 32'h576439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2932   :   assert (rdbk == 32'hccca7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2933   :   assert (rdbk == 32'h525a2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2934   :   assert (rdbk == 32'h5cb98d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2935   :   assert (rdbk == 32'h7dd99f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2936   :   assert (rdbk == 32'h164b85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2937   :   assert (rdbk == 32'h28a0b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2938   :   assert (rdbk == 32'h73c5a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2939   :   assert (rdbk == 32'h496daa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2940   :   assert (rdbk == 32'h3b991d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2941   :   assert (rdbk == 32'h35b6a1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2942   :   assert (rdbk == 32'h2d429d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2943   :   assert (rdbk == 32'h250318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2944   :   assert (rdbk == 32'h7c1ffe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2945   :   assert (rdbk == 32'h27c29e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2946   :   assert (rdbk == 32'h79eda2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2947   :   assert (rdbk == 32'h70fc3f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2948   :   assert (rdbk == 32'h56be63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2949   :   assert (rdbk == 32'h625671) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2950   :   assert (rdbk == 32'h5d3c56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2951   :   assert (rdbk == 32'h10cabc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2952   :   assert (rdbk == 32'h526336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2953   :   assert (rdbk == 32'h167737) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2954   :   assert (rdbk == 32'h2f3cd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2955   :   assert (rdbk == 32'h2884e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2956   :   assert (rdbk == 32'h779f64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2957   :   assert (rdbk == 32'h2002e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2958   :   assert (rdbk == 32'h5dd9f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2959   :   assert (rdbk == 32'h578c30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2960   :   assert (rdbk == 32'h4fe90e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2961   :   assert (rdbk == 32'h5dd571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2962   :   assert (rdbk == 32'h1efe54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2963   :   assert (rdbk == 32'h3b819b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2964   :   assert (rdbk == 32'h55cf42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2965   :   assert (rdbk == 32'h7c6280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2966   :   assert (rdbk == 32'h4c16a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2967   :   assert (rdbk == 32'h681118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2968   :   assert (rdbk == 32'h3512d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2969   :   assert (rdbk == 32'h48464d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2970   :   assert (rdbk == 32'h58ba3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2971   :   assert (rdbk == 32'h5d5408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2972   :   assert (rdbk == 32'h6d8c9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2973   :   assert (rdbk == 32'h60f339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2974   :   assert (rdbk == 32'h472ec9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2975   :   assert (rdbk == 32'h6b65a9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2976   :   assert (rdbk == 32'h72084b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2977   :   assert (rdbk == 32'h5a063f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2978   :   assert (rdbk == 32'h43655b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2979   :   assert (rdbk == 32'h6e099c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2980   :   assert (rdbk == 32'h66cfc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2981   :   assert (rdbk == 32'h3a288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2982   :   assert (rdbk == 32'he8f2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2983   :   assert (rdbk == 32'h5fe774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2984   :   assert (rdbk == 32'h5532aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2985   :   assert (rdbk == 32'h1eb08a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2986   :   assert (rdbk == 32'h72b2c6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2987   :   assert (rdbk == 32'h3680d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2988   :   assert (rdbk == 32'h35fe5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2989   :   assert (rdbk == 32'h6fc477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2990   :   assert (rdbk == 32'h7b9d9f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2991   :   assert (rdbk == 32'h479572) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2992   :   assert (rdbk == 32'h36b40e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2993   :   assert (rdbk == 32'h45d67a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2994   :   assert (rdbk == 32'h3e8ae1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2995   :   assert (rdbk == 32'h79f13d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2996   :   assert (rdbk == 32'h1eed4d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2997   :   assert (rdbk == 32'h4a65e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2998   :   assert (rdbk == 32'h1fc634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	2999   :   assert (rdbk == 32'h20a59f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3000   :   assert (rdbk == 32'h777efb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3001   :   assert (rdbk == 32'h2ac58c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3002   :   assert (rdbk == 32'h33c85e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3003   :   assert (rdbk == 32'h57c20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3004   :   assert (rdbk == 32'h72f8ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3005   :   assert (rdbk == 32'he1477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3006   :   assert (rdbk == 32'h314108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3007   :   assert (rdbk == 32'h2792bb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3008   :   assert (rdbk == 32'h43ebcb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3009   :   assert (rdbk == 32'h3174aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3010   :   assert (rdbk == 32'h24e42f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3011   :   assert (rdbk == 32'h4b8aaf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3012   :   assert (rdbk == 32'h4a971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3013   :   assert (rdbk == 32'h18bff5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3014   :   assert (rdbk == 32'h3fcafa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3015   :   assert (rdbk == 32'h32ee93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3016   :   assert (rdbk == 32'h6c6b5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3017   :   assert (rdbk == 32'h3f20a9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3018   :   assert (rdbk == 32'h2f666c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3019   :   assert (rdbk == 32'h59a287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3020   :   assert (rdbk == 32'h3c4941) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3021   :   assert (rdbk == 32'h6fecec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3022   :   assert (rdbk == 32'h3ed865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3023   :   assert (rdbk == 32'h1fa265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3024   :   assert (rdbk == 32'h19c27f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3025   :   assert (rdbk == 32'h49e8e1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3026   :   assert (rdbk == 32'h11c03b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3027   :   assert (rdbk == 32'h7c669f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3028   :   assert (rdbk == 32'h4dae9d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3029   :   assert (rdbk == 32'h5a457f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3030   :   assert (rdbk == 32'h6072) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3031   :   assert (rdbk == 32'h308862) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3032   :   assert (rdbk == 32'h67b6a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3033   :   assert (rdbk == 32'h55b1d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3034   :   assert (rdbk == 32'h6e642f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3035   :   assert (rdbk == 32'h1da8e2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3036   :   assert (rdbk == 32'h4aad61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3037   :   assert (rdbk == 32'h7ba2d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3038   :   assert (rdbk == 32'h22becf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3039   :   assert (rdbk == 32'h89007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3040   :   assert (rdbk == 32'h24159d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3041   :   assert (rdbk == 32'h118c4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3042   :   assert (rdbk == 32'h49fcd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3043   :   assert (rdbk == 32'h7cd6f8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3044   :   assert (rdbk == 32'hee1ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3045   :   assert (rdbk == 32'h343c50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3046   :   assert (rdbk == 32'h5e6088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3047   :   assert (rdbk == 32'h39cb93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3048   :   assert (rdbk == 32'h4442da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3049   :   assert (rdbk == 32'h5633df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3050   :   assert (rdbk == 32'h6cb923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3051   :   assert (rdbk == 32'h39b6b1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3052   :   assert (rdbk == 32'h15ed43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3053   :   assert (rdbk == 32'h5e7e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3054   :   assert (rdbk == 32'h6920a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3055   :   assert (rdbk == 32'h2637df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3056   :   assert (rdbk == 32'h4040da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3057   :   assert (rdbk == 32'h6a4bea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3058   :   assert (rdbk == 32'h4fda40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3059   :   assert (rdbk == 32'h50aa86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3060   :   assert (rdbk == 32'h587b50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3061   :   assert (rdbk == 32'h770c2d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3062   :   assert (rdbk == 32'h198a5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3063   :   assert (rdbk == 32'h484497) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3064   :   assert (rdbk == 32'h26c491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3065   :   assert (rdbk == 32'h31f27b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3066   :   assert (rdbk == 32'h661e20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3067   :   assert (rdbk == 32'h497637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3068   :   assert (rdbk == 32'h3e64cd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3069   :   assert (rdbk == 32'h11644d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3070   :   assert (rdbk == 32'h4dbf5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3071   :   assert (rdbk == 32'h5d3b5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h300
	3072   :   assert (rdbk == 32'h54ba24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3073   :   assert (rdbk == 32'h105da7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3074   :   assert (rdbk == 32'h1820c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3075   :   assert (rdbk == 32'h563458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3076   :   assert (rdbk == 32'h182c86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3077   :   assert (rdbk == 32'h5a9e87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3078   :   assert (rdbk == 32'h2b3243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3079   :   assert (rdbk == 32'h7d6401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3080   :   assert (rdbk == 32'h380bfc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3081   :   assert (rdbk == 32'h4642b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3082   :   assert (rdbk == 32'h6a49f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3083   :   assert (rdbk == 32'h71c01d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3084   :   assert (rdbk == 32'h7c54cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3085   :   assert (rdbk == 32'h6a447c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3086   :   assert (rdbk == 32'h733a13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3087   :   assert (rdbk == 32'h1ff309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3088   :   assert (rdbk == 32'h17637c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3089   :   assert (rdbk == 32'h403603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3090   :   assert (rdbk == 32'hd378f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3091   :   assert (rdbk == 32'h502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3092   :   assert (rdbk == 32'h78738f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3093   :   assert (rdbk == 32'h2d3acc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3094   :   assert (rdbk == 32'h4c9458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3095   :   assert (rdbk == 32'h26636f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3096   :   assert (rdbk == 32'h4fb661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3097   :   assert (rdbk == 32'h4300ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3098   :   assert (rdbk == 32'h205f41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3099   :   assert (rdbk == 32'h1fde13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3100   :   assert (rdbk == 32'h2a5d85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3101   :   assert (rdbk == 32'h78f33e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3102   :   assert (rdbk == 32'hd9202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3103   :   assert (rdbk == 32'h2e81bf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3104   :   assert (rdbk == 32'h1bcc4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3105   :   assert (rdbk == 32'h2cd5ad) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3106   :   assert (rdbk == 32'h115ddf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3107   :   assert (rdbk == 32'h4aa7ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3108   :   assert (rdbk == 32'h26734f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3109   :   assert (rdbk == 32'h574417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3110   :   assert (rdbk == 32'h697d18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3111   :   assert (rdbk == 32'h70a8ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3112   :   assert (rdbk == 32'h7cb0eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3113   :   assert (rdbk == 32'h1e94c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3114   :   assert (rdbk == 32'h7f89d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3115   :   assert (rdbk == 32'h1129fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3116   :   assert (rdbk == 32'h5b1e76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3117   :   assert (rdbk == 32'h6c0abc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3118   :   assert (rdbk == 32'h17b7ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3119   :   assert (rdbk == 32'h67992c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3120   :   assert (rdbk == 32'h3df38a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3121   :   assert (rdbk == 32'h7af33f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3122   :   assert (rdbk == 32'hfb6a9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3123   :   assert (rdbk == 32'h43a165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3124   :   assert (rdbk == 32'h37e04) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3125   :   assert (rdbk == 32'h172ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3126   :   assert (rdbk == 32'h3e29a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3127   :   assert (rdbk == 32'h1bc9fe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3128   :   assert (rdbk == 32'h3e135f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3129   :   assert (rdbk == 32'h6a9b05) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3130   :   assert (rdbk == 32'h55a9db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3131   :   assert (rdbk == 32'h30ebbb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3132   :   assert (rdbk == 32'h2fc89a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3133   :   assert (rdbk == 32'h1e3dea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3134   :   assert (rdbk == 32'h76426c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3135   :   assert (rdbk == 32'h26893b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3136   :   assert (rdbk == 32'h3f2681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3137   :   assert (rdbk == 32'h63c7ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3138   :   assert (rdbk == 32'he7b22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3139   :   assert (rdbk == 32'h86a72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3140   :   assert (rdbk == 32'h466061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3141   :   assert (rdbk == 32'h661226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3142   :   assert (rdbk == 32'h244178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3143   :   assert (rdbk == 32'h4d8373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3144   :   assert (rdbk == 32'h6ae00e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3145   :   assert (rdbk == 32'h437707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3146   :   assert (rdbk == 32'h1f1551) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3147   :   assert (rdbk == 32'h209652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3148   :   assert (rdbk == 32'h5aba83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3149   :   assert (rdbk == 32'h35e5b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3150   :   assert (rdbk == 32'h50c34f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3151   :   assert (rdbk == 32'h3dcc54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3152   :   assert (rdbk == 32'h51e1a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3153   :   assert (rdbk == 32'h44755a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3154   :   assert (rdbk == 32'h502ed5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3155   :   assert (rdbk == 32'h7f0280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3156   :   assert (rdbk == 32'h100f23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3157   :   assert (rdbk == 32'h2ffa94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3158   :   assert (rdbk == 32'h1d1ade) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3159   :   assert (rdbk == 32'h4a5b7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3160   :   assert (rdbk == 32'h14c483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3161   :   assert (rdbk == 32'h197f8c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3162   :   assert (rdbk == 32'h68dfdc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3163   :   assert (rdbk == 32'h39c644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3164   :   assert (rdbk == 32'h213e7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3165   :   assert (rdbk == 32'h20cfce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3166   :   assert (rdbk == 32'h69a2a1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3167   :   assert (rdbk == 32'h5dcd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3168   :   assert (rdbk == 32'h9f2cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3169   :   assert (rdbk == 32'h59a23b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3170   :   assert (rdbk == 32'h737888) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3171   :   assert (rdbk == 32'h56886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3172   :   assert (rdbk == 32'h55ca97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3173   :   assert (rdbk == 32'h3a3788) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3174   :   assert (rdbk == 32'h7dc26e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3175   :   assert (rdbk == 32'h7e3dfe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3176   :   assert (rdbk == 32'h3a2d39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3177   :   assert (rdbk == 32'h318c68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3178   :   assert (rdbk == 32'h5a687e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3179   :   assert (rdbk == 32'h38c275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3180   :   assert (rdbk == 32'h38decf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3181   :   assert (rdbk == 32'h2f9c8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3182   :   assert (rdbk == 32'h254843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3183   :   assert (rdbk == 32'h5084b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3184   :   assert (rdbk == 32'h4c8908) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3185   :   assert (rdbk == 32'h58b784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3186   :   assert (rdbk == 32'h413c8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3187   :   assert (rdbk == 32'he6e75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3188   :   assert (rdbk == 32'h455752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3189   :   assert (rdbk == 32'h12af11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3190   :   assert (rdbk == 32'h2669c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3191   :   assert (rdbk == 32'h5172c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3192   :   assert (rdbk == 32'h2215d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3193   :   assert (rdbk == 32'h2819df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3194   :   assert (rdbk == 32'h786948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3195   :   assert (rdbk == 32'h606a08) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3196   :   assert (rdbk == 32'h22c575) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3197   :   assert (rdbk == 32'h5bfc40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3198   :   assert (rdbk == 32'h103084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3199   :   assert (rdbk == 32'h546138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3200   :   assert (rdbk == 32'h45c01c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3201   :   assert (rdbk == 32'h7302e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3202   :   assert (rdbk == 32'h2c486c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3203   :   assert (rdbk == 32'h566959) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3204   :   assert (rdbk == 32'h75417e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3205   :   assert (rdbk == 32'h45b76e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3206   :   assert (rdbk == 32'h7977af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3207   :   assert (rdbk == 32'h513803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3208   :   assert (rdbk == 32'h39bef8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3209   :   assert (rdbk == 32'h4b900e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3210   :   assert (rdbk == 32'h46d2fc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3211   :   assert (rdbk == 32'h400a68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3212   :   assert (rdbk == 32'h4d6515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3213   :   assert (rdbk == 32'h78e1e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3214   :   assert (rdbk == 32'h44ef74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3215   :   assert (rdbk == 32'h327a8d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3216   :   assert (rdbk == 32'h31f23d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3217   :   assert (rdbk == 32'h62c1ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3218   :   assert (rdbk == 32'h1c6133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3219   :   assert (rdbk == 32'h683de5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3220   :   assert (rdbk == 32'h501b1f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3221   :   assert (rdbk == 32'h52a8a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3222   :   assert (rdbk == 32'h267789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3223   :   assert (rdbk == 32'h415d50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3224   :   assert (rdbk == 32'h8abab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3225   :   assert (rdbk == 32'h1e6b4f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3226   :   assert (rdbk == 32'h6a8345) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3227   :   assert (rdbk == 32'h47d3f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3228   :   assert (rdbk == 32'h6fe5cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3229   :   assert (rdbk == 32'h6e826b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3230   :   assert (rdbk == 32'h193852) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3231   :   assert (rdbk == 32'h89a79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3232   :   assert (rdbk == 32'h2bb422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3233   :   assert (rdbk == 32'h126a56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3234   :   assert (rdbk == 32'h7be58c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3235   :   assert (rdbk == 32'h43e2a4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3236   :   assert (rdbk == 32'hf8b38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3237   :   assert (rdbk == 32'h1b2b4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3238   :   assert (rdbk == 32'h2c667f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3239   :   assert (rdbk == 32'ha45dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3240   :   assert (rdbk == 32'h56743f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3241   :   assert (rdbk == 32'h1ead18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3242   :   assert (rdbk == 32'h7a2b5e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3243   :   assert (rdbk == 32'h76bd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3244   :   assert (rdbk == 32'h2a3bee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3245   :   assert (rdbk == 32'h590a3d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3246   :   assert (rdbk == 32'h71bcf2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3247   :   assert (rdbk == 32'h18eadb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3248   :   assert (rdbk == 32'h1eaefb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3249   :   assert (rdbk == 32'h4aec0f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3250   :   assert (rdbk == 32'h3208d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3251   :   assert (rdbk == 32'h361f53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3252   :   assert (rdbk == 32'h18c89a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3253   :   assert (rdbk == 32'h2664db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3254   :   assert (rdbk == 32'h4f52e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3255   :   assert (rdbk == 32'h27ba5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3256   :   assert (rdbk == 32'h6333ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3257   :   assert (rdbk == 32'hf088b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3258   :   assert (rdbk == 32'h2d6fbc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3259   :   assert (rdbk == 32'h75acd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3260   :   assert (rdbk == 32'h74d672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3261   :   assert (rdbk == 32'h6d4d35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3262   :   assert (rdbk == 32'h9188c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3263   :   assert (rdbk == 32'h7d5aa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3264   :   assert (rdbk == 32'h1ef3df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3265   :   assert (rdbk == 32'h1f9af3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3266   :   assert (rdbk == 32'h10535e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3267   :   assert (rdbk == 32'h7e31cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3268   :   assert (rdbk == 32'h77dec7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3269   :   assert (rdbk == 32'h6e71a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3270   :   assert (rdbk == 32'h781b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3271   :   assert (rdbk == 32'h4b4ce5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3272   :   assert (rdbk == 32'h20d5ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3273   :   assert (rdbk == 32'h38b2f9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3274   :   assert (rdbk == 32'h48c010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3275   :   assert (rdbk == 32'h122894) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3276   :   assert (rdbk == 32'h72fed3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3277   :   assert (rdbk == 32'h717ddb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3278   :   assert (rdbk == 32'h646008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3279   :   assert (rdbk == 32'h374436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3280   :   assert (rdbk == 32'h7e60b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3281   :   assert (rdbk == 32'h4d7b55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3282   :   assert (rdbk == 32'h95348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3283   :   assert (rdbk == 32'h1ef29e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3284   :   assert (rdbk == 32'h542939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3285   :   assert (rdbk == 32'hb916a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3286   :   assert (rdbk == 32'h290ffa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3287   :   assert (rdbk == 32'h48f557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3288   :   assert (rdbk == 32'h3c0a36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3289   :   assert (rdbk == 32'h141f7e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3290   :   assert (rdbk == 32'h3dbaac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3291   :   assert (rdbk == 32'h3abfa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3292   :   assert (rdbk == 32'h7db465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3293   :   assert (rdbk == 32'h3dfe71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3294   :   assert (rdbk == 32'h130ac5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3295   :   assert (rdbk == 32'h66c748) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3296   :   assert (rdbk == 32'h439d62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3297   :   assert (rdbk == 32'h70a8ce) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3298   :   assert (rdbk == 32'h6e41a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3299   :   assert (rdbk == 32'h4b1959) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3300   :   assert (rdbk == 32'h689661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3301   :   assert (rdbk == 32'h793677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3302   :   assert (rdbk == 32'h265e13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3303   :   assert (rdbk == 32'h2dbac6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3304   :   assert (rdbk == 32'h42f829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3305   :   assert (rdbk == 32'h20829c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3306   :   assert (rdbk == 32'h510f7b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3307   :   assert (rdbk == 32'h4ec4fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3308   :   assert (rdbk == 32'h25509c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3309   :   assert (rdbk == 32'h43b57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3310   :   assert (rdbk == 32'h5aa08f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3311   :   assert (rdbk == 32'h6a3cb4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3312   :   assert (rdbk == 32'h26578b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3313   :   assert (rdbk == 32'h759ee8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3314   :   assert (rdbk == 32'h20f02f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3315   :   assert (rdbk == 32'h30256c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3316   :   assert (rdbk == 32'h76ebb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3317   :   assert (rdbk == 32'h7df826) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3318   :   assert (rdbk == 32'h6d0719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3319   :   assert (rdbk == 32'h6e712e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3320   :   assert (rdbk == 32'h390d6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3321   :   assert (rdbk == 32'h76cf37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3322   :   assert (rdbk == 32'h58e4b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3323   :   assert (rdbk == 32'h1a0d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3324   :   assert (rdbk == 32'h323629) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3325   :   assert (rdbk == 32'h269540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3326   :   assert (rdbk == 32'h29787a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3327   :   assert (rdbk == 32'h2ac3e4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h301
	3328   :   assert (rdbk == 32'hbd73b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3329   :   assert (rdbk == 32'h6e6ff2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3330   :   assert (rdbk == 32'h33b73d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3331   :   assert (rdbk == 32'h18142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3332   :   assert (rdbk == 32'h37c055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3333   :   assert (rdbk == 32'hc793a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3334   :   assert (rdbk == 32'h63d54c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3335   :   assert (rdbk == 32'h65b53b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3336   :   assert (rdbk == 32'h2b6d22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3337   :   assert (rdbk == 32'h276756) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3338   :   assert (rdbk == 32'hbf850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3339   :   assert (rdbk == 32'h371eb7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3340   :   assert (rdbk == 32'h7e0eae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3341   :   assert (rdbk == 32'h55f447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3342   :   assert (rdbk == 32'h2c6478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3343   :   assert (rdbk == 32'h762f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3344   :   assert (rdbk == 32'h1954f8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3345   :   assert (rdbk == 32'h2aceeb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3346   :   assert (rdbk == 32'h5a8c95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3347   :   assert (rdbk == 32'h59c893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3348   :   assert (rdbk == 32'h7ad993) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3349   :   assert (rdbk == 32'h3fcc6b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3350   :   assert (rdbk == 32'h3bb28d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3351   :   assert (rdbk == 32'h17c70b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3352   :   assert (rdbk == 32'h3472d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3353   :   assert (rdbk == 32'h524746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3354   :   assert (rdbk == 32'h3d5aa2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3355   :   assert (rdbk == 32'h496fd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3356   :   assert (rdbk == 32'h2ce2fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3357   :   assert (rdbk == 32'h7b9b75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3358   :   assert (rdbk == 32'h645e08) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3359   :   assert (rdbk == 32'h271c00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3360   :   assert (rdbk == 32'h5f5790) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3361   :   assert (rdbk == 32'h1d6259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3362   :   assert (rdbk == 32'h61845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3363   :   assert (rdbk == 32'h58b886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3364   :   assert (rdbk == 32'h667d07) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3365   :   assert (rdbk == 32'h2e64e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3366   :   assert (rdbk == 32'h7a6345) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3367   :   assert (rdbk == 32'h603ef6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3368   :   assert (rdbk == 32'h3ca9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3369   :   assert (rdbk == 32'h4ae8b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3370   :   assert (rdbk == 32'h364ffa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3371   :   assert (rdbk == 32'h773af1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3372   :   assert (rdbk == 32'h5d1dcf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3373   :   assert (rdbk == 32'h75525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3374   :   assert (rdbk == 32'h3d2500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3375   :   assert (rdbk == 32'h660416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3376   :   assert (rdbk == 32'h39905c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3377   :   assert (rdbk == 32'h7921f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3378   :   assert (rdbk == 32'h3e43ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3379   :   assert (rdbk == 32'h60b05f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3380   :   assert (rdbk == 32'h4f50c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3381   :   assert (rdbk == 32'h2f3124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3382   :   assert (rdbk == 32'h3546ed) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3383   :   assert (rdbk == 32'h77a145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3384   :   assert (rdbk == 32'h6fe39f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3385   :   assert (rdbk == 32'h76fbfc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3386   :   assert (rdbk == 32'h649e75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3387   :   assert (rdbk == 32'h640f8e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3388   :   assert (rdbk == 32'h1bbb26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3389   :   assert (rdbk == 32'h5c1abd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3390   :   assert (rdbk == 32'h172189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3391   :   assert (rdbk == 32'h19bc1f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3392   :   assert (rdbk == 32'h419408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3393   :   assert (rdbk == 32'h7a08cb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3394   :   assert (rdbk == 32'h6d03f9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3395   :   assert (rdbk == 32'h5c228d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3396   :   assert (rdbk == 32'h62ded2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3397   :   assert (rdbk == 32'h3799af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3398   :   assert (rdbk == 32'h362d26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3399   :   assert (rdbk == 32'h189939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3400   :   assert (rdbk == 32'h4d7c96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3401   :   assert (rdbk == 32'hf2040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3402   :   assert (rdbk == 32'h24a232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3403   :   assert (rdbk == 32'h710d5d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3404   :   assert (rdbk == 32'h326c77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3405   :   assert (rdbk == 32'h346c07) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3406   :   assert (rdbk == 32'h3b6d44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3407   :   assert (rdbk == 32'h6312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3408   :   assert (rdbk == 32'h3fa9a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3409   :   assert (rdbk == 32'h582478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3410   :   assert (rdbk == 32'h7df703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3411   :   assert (rdbk == 32'h682c9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3412   :   assert (rdbk == 32'h339be2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3413   :   assert (rdbk == 32'h799c05) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3414   :   assert (rdbk == 32'h12b0b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3415   :   assert (rdbk == 32'h57bbe) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3416   :   assert (rdbk == 32'h3b85e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3417   :   assert (rdbk == 32'h2d1369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3418   :   assert (rdbk == 32'h7cc14c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3419   :   assert (rdbk == 32'h78df50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3420   :   assert (rdbk == 32'h42dc00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3421   :   assert (rdbk == 32'h38605c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3422   :   assert (rdbk == 32'h4e1b34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3423   :   assert (rdbk == 32'h13a1a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3424   :   assert (rdbk == 32'h6c1a74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3425   :   assert (rdbk == 32'h10a618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3426   :   assert (rdbk == 32'h2c96ae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3427   :   assert (rdbk == 32'h7e9d89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3428   :   assert (rdbk == 32'h371ac9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3429   :   assert (rdbk == 32'h3c6b6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3430   :   assert (rdbk == 32'h22b503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3431   :   assert (rdbk == 32'h14e72b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3432   :   assert (rdbk == 32'h2de608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3433   :   assert (rdbk == 32'hce903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3434   :   assert (rdbk == 32'h5d40d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3435   :   assert (rdbk == 32'hdce8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3436   :   assert (rdbk == 32'h18b97a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3437   :   assert (rdbk == 32'he2866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3438   :   assert (rdbk == 32'h25bb61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3439   :   assert (rdbk == 32'h4e7810) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3440   :   assert (rdbk == 32'h268c8c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3441   :   assert (rdbk == 32'h12bf94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3442   :   assert (rdbk == 32'h34678c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3443   :   assert (rdbk == 32'h38b9e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3444   :   assert (rdbk == 32'h18b648) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3445   :   assert (rdbk == 32'h55917c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3446   :   assert (rdbk == 32'h6f6840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3447   :   assert (rdbk == 32'h30ad0e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3448   :   assert (rdbk == 32'h5f32ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3449   :   assert (rdbk == 32'h67e44e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3450   :   assert (rdbk == 32'h372d52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3451   :   assert (rdbk == 32'hd8f9a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3452   :   assert (rdbk == 32'h32d614) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3453   :   assert (rdbk == 32'h282e2f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3454   :   assert (rdbk == 32'h51b18a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3455   :   assert (rdbk == 32'h3be2ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3456   :   assert (rdbk == 32'h45e1a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3457   :   assert (rdbk == 32'h4f9a0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3458   :   assert (rdbk == 32'h304cc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3459   :   assert (rdbk == 32'h45f4c2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3460   :   assert (rdbk == 32'h15ad78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3461   :   assert (rdbk == 32'h20c3f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3462   :   assert (rdbk == 32'h6d7b58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3463   :   assert (rdbk == 32'hcb84e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3464   :   assert (rdbk == 32'h35214e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3465   :   assert (rdbk == 32'h179161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3466   :   assert (rdbk == 32'h3fd456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3467   :   assert (rdbk == 32'h7dac64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3468   :   assert (rdbk == 32'h5c65ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3469   :   assert (rdbk == 32'h462b00) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3470   :   assert (rdbk == 32'h265667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3471   :   assert (rdbk == 32'h6d98a9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3472   :   assert (rdbk == 32'h41c118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3473   :   assert (rdbk == 32'h5b3c27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3474   :   assert (rdbk == 32'h6ad6fd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3475   :   assert (rdbk == 32'h1cdf1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3476   :   assert (rdbk == 32'h163f26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3477   :   assert (rdbk == 32'h424ec7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3478   :   assert (rdbk == 32'h475985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3479   :   assert (rdbk == 32'h13acba) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3480   :   assert (rdbk == 32'h662217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3481   :   assert (rdbk == 32'h566c12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3482   :   assert (rdbk == 32'h63afe6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3483   :   assert (rdbk == 32'h5e3106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3484   :   assert (rdbk == 32'h4f0daa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3485   :   assert (rdbk == 32'h46e674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3486   :   assert (rdbk == 32'h7d366d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3487   :   assert (rdbk == 32'h57917d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3488   :   assert (rdbk == 32'h63c474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3489   :   assert (rdbk == 32'h1056a2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3490   :   assert (rdbk == 32'h79be96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3491   :   assert (rdbk == 32'h25de7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3492   :   assert (rdbk == 32'h50d646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3493   :   assert (rdbk == 32'h58c72c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3494   :   assert (rdbk == 32'h32e26b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3495   :   assert (rdbk == 32'h600242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3496   :   assert (rdbk == 32'h1c5fae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3497   :   assert (rdbk == 32'h4894bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3498   :   assert (rdbk == 32'h136910) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3499   :   assert (rdbk == 32'h41d11a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3500   :   assert (rdbk == 32'h3a6309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3501   :   assert (rdbk == 32'h339bb0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3502   :   assert (rdbk == 32'h509990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3503   :   assert (rdbk == 32'h69ae48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3504   :   assert (rdbk == 32'h3dbd23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3505   :   assert (rdbk == 32'h3c2459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3506   :   assert (rdbk == 32'h7c0511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3507   :   assert (rdbk == 32'h1fca94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3508   :   assert (rdbk == 32'h6ac48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3509   :   assert (rdbk == 32'h7cd3e1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3510   :   assert (rdbk == 32'h60b8bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3511   :   assert (rdbk == 32'h53ce37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3512   :   assert (rdbk == 32'h770423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3513   :   assert (rdbk == 32'h187742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3514   :   assert (rdbk == 32'h77a150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3515   :   assert (rdbk == 32'h2b0b33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3516   :   assert (rdbk == 32'h61b6fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3517   :   assert (rdbk == 32'h573ef8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3518   :   assert (rdbk == 32'h547fff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3519   :   assert (rdbk == 32'h1f486e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3520   :   assert (rdbk == 32'h7dd70a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3521   :   assert (rdbk == 32'h378642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3522   :   assert (rdbk == 32'h34e5f8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3523   :   assert (rdbk == 32'h27d2df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3524   :   assert (rdbk == 32'h58a86c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3525   :   assert (rdbk == 32'h63153d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3526   :   assert (rdbk == 32'h2f742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3527   :   assert (rdbk == 32'h267dae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3528   :   assert (rdbk == 32'h330b1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3529   :   assert (rdbk == 32'h3cdc41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3530   :   assert (rdbk == 32'h46cd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3531   :   assert (rdbk == 32'h2f61c4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3532   :   assert (rdbk == 32'h6b68f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3533   :   assert (rdbk == 32'h2f18c8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3534   :   assert (rdbk == 32'h5e02ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3535   :   assert (rdbk == 32'h5d25cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3536   :   assert (rdbk == 32'h1d0fd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3537   :   assert (rdbk == 32'h611371) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3538   :   assert (rdbk == 32'h6c6620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3539   :   assert (rdbk == 32'h6e786e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3540   :   assert (rdbk == 32'h44c168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3541   :   assert (rdbk == 32'h74c99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3542   :   assert (rdbk == 32'h6d81e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3543   :   assert (rdbk == 32'hef14e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3544   :   assert (rdbk == 32'h7dc101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3545   :   assert (rdbk == 32'h65e2e0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3546   :   assert (rdbk == 32'h5f8a06) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3547   :   assert (rdbk == 32'h566e0a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3548   :   assert (rdbk == 32'h46e620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3549   :   assert (rdbk == 32'h21a654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3550   :   assert (rdbk == 32'h23c537) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3551   :   assert (rdbk == 32'h57bb45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3552   :   assert (rdbk == 32'h3136e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3553   :   assert (rdbk == 32'h1cb61a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3554   :   assert (rdbk == 32'h606f86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3555   :   assert (rdbk == 32'h1ef140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3556   :   assert (rdbk == 32'h5b911d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3557   :   assert (rdbk == 32'h32970f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3558   :   assert (rdbk == 32'h5f2593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3559   :   assert (rdbk == 32'h3932f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3560   :   assert (rdbk == 32'h34020f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3561   :   assert (rdbk == 32'hdbbea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3562   :   assert (rdbk == 32'h46615c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3563   :   assert (rdbk == 32'h15a1e9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3564   :   assert (rdbk == 32'h1b005d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3565   :   assert (rdbk == 32'h1df31a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3566   :   assert (rdbk == 32'h604ae9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3567   :   assert (rdbk == 32'h1f8d6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3568   :   assert (rdbk == 32'h594dc1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3569   :   assert (rdbk == 32'h2c0e16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3570   :   assert (rdbk == 32'h32bff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3571   :   assert (rdbk == 32'h588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3572   :   assert (rdbk == 32'h1b614d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3573   :   assert (rdbk == 32'h4a7d11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3574   :   assert (rdbk == 32'h33b785) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3575   :   assert (rdbk == 32'h63c1e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3576   :   assert (rdbk == 32'h585159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3577   :   assert (rdbk == 32'h75da02) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3578   :   assert (rdbk == 32'h43fad0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3579   :   assert (rdbk == 32'h180399) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3580   :   assert (rdbk == 32'h7dc9f9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3581   :   assert (rdbk == 32'h3fbb7a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3582   :   assert (rdbk == 32'h7d233b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3583   :   assert (rdbk == 32'h6c4e15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h302
	3584   :   assert (rdbk == 32'h7528df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3585   :   assert (rdbk == 32'h27e542) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3586   :   assert (rdbk == 32'h61ae1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3587   :   assert (rdbk == 32'he7619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3588   :   assert (rdbk == 32'h2a2121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3589   :   assert (rdbk == 32'h6e8b13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3590   :   assert (rdbk == 32'h680dfa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3591   :   assert (rdbk == 32'h40e4db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3592   :   assert (rdbk == 32'h34b45f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3593   :   assert (rdbk == 32'h11f605) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3594   :   assert (rdbk == 32'h46f89d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3595   :   assert (rdbk == 32'h1e81af) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3596   :   assert (rdbk == 32'h4a250c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3597   :   assert (rdbk == 32'h7b37cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3598   :   assert (rdbk == 32'h71ec72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3599   :   assert (rdbk == 32'h4394b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3600   :   assert (rdbk == 32'h66bee0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3601   :   assert (rdbk == 32'h56fa73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3602   :   assert (rdbk == 32'h7a2ea3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3603   :   assert (rdbk == 32'h533298) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3604   :   assert (rdbk == 32'h631199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3605   :   assert (rdbk == 32'h3e3c7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3606   :   assert (rdbk == 32'h3cc584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3607   :   assert (rdbk == 32'h490773) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3608   :   assert (rdbk == 32'h2cbd2b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3609   :   assert (rdbk == 32'h40dc2e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3610   :   assert (rdbk == 32'h300f57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3611   :   assert (rdbk == 32'h21fffc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3612   :   assert (rdbk == 32'h3a9a09) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3613   :   assert (rdbk == 32'h1d90e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3614   :   assert (rdbk == 32'h4d017b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3615   :   assert (rdbk == 32'h4e9991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3616   :   assert (rdbk == 32'h64b2ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3617   :   assert (rdbk == 32'h5ab4f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3618   :   assert (rdbk == 32'hf271c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3619   :   assert (rdbk == 32'h30e7b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3620   :   assert (rdbk == 32'h4fd31e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3621   :   assert (rdbk == 32'h5c4d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3622   :   assert (rdbk == 32'h221801) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3623   :   assert (rdbk == 32'h425e76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3624   :   assert (rdbk == 32'h47d7ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3625   :   assert (rdbk == 32'h18b679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3626   :   assert (rdbk == 32'he3bbf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3627   :   assert (rdbk == 32'h14166c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3628   :   assert (rdbk == 32'h125f1a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3629   :   assert (rdbk == 32'h624156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3630   :   assert (rdbk == 32'h58b498) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3631   :   assert (rdbk == 32'h77f737) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3632   :   assert (rdbk == 32'hde09e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3633   :   assert (rdbk == 32'h5a1403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3634   :   assert (rdbk == 32'h22dd7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3635   :   assert (rdbk == 32'h6d51a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3636   :   assert (rdbk == 32'h4a18a0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3637   :   assert (rdbk == 32'hd9bb9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3638   :   assert (rdbk == 32'h59d1b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3639   :   assert (rdbk == 32'h14ab6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3640   :   assert (rdbk == 32'h75264d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3641   :   assert (rdbk == 32'h5fed95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3642   :   assert (rdbk == 32'h50fb2f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3643   :   assert (rdbk == 32'h3fd33d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3644   :   assert (rdbk == 32'h7af46c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3645   :   assert (rdbk == 32'h33315f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3646   :   assert (rdbk == 32'h5adbcc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3647   :   assert (rdbk == 32'h78e07) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3648   :   assert (rdbk == 32'h64e37d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3649   :   assert (rdbk == 32'h324918) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3650   :   assert (rdbk == 32'h7caa8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3651   :   assert (rdbk == 32'h28ed0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3652   :   assert (rdbk == 32'h2b84bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3653   :   assert (rdbk == 32'h500889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3654   :   assert (rdbk == 32'h2fba24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3655   :   assert (rdbk == 32'h4dfd0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3656   :   assert (rdbk == 32'h41b5c6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3657   :   assert (rdbk == 32'h4330a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3658   :   assert (rdbk == 32'h41c081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3659   :   assert (rdbk == 32'h3f3704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3660   :   assert (rdbk == 32'h7e234d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3661   :   assert (rdbk == 32'h795a1a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3662   :   assert (rdbk == 32'h4ed76c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3663   :   assert (rdbk == 32'h8ad40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3664   :   assert (rdbk == 32'h4d4d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3665   :   assert (rdbk == 32'h98c2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3666   :   assert (rdbk == 32'h2c462d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3667   :   assert (rdbk == 32'h7d999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3668   :   assert (rdbk == 32'h2e6131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3669   :   assert (rdbk == 32'h6ebf5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3670   :   assert (rdbk == 32'h555cf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3671   :   assert (rdbk == 32'h34f5df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3672   :   assert (rdbk == 32'h7ed5c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3673   :   assert (rdbk == 32'h3871b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3674   :   assert (rdbk == 32'h9f9d8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3675   :   assert (rdbk == 32'h21816b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3676   :   assert (rdbk == 32'h996e1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3677   :   assert (rdbk == 32'h29874c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3678   :   assert (rdbk == 32'h6f4069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3679   :   assert (rdbk == 32'h521ae5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3680   :   assert (rdbk == 32'h2419f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3681   :   assert (rdbk == 32'h4bb714) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3682   :   assert (rdbk == 32'h230e90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3683   :   assert (rdbk == 32'h372eb3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3684   :   assert (rdbk == 32'h3c737c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3685   :   assert (rdbk == 32'h5ad44b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3686   :   assert (rdbk == 32'h64f614) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3687   :   assert (rdbk == 32'h3ed2d1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3688   :   assert (rdbk == 32'h143636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3689   :   assert (rdbk == 32'h4b8d3d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3690   :   assert (rdbk == 32'h78bf78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3691   :   assert (rdbk == 32'h87600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3692   :   assert (rdbk == 32'h12f761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3693   :   assert (rdbk == 32'h54fd7c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3694   :   assert (rdbk == 32'hd02de) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3695   :   assert (rdbk == 32'h50ad17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3696   :   assert (rdbk == 32'h44930c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3697   :   assert (rdbk == 32'h671632) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3698   :   assert (rdbk == 32'h1360bd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3699   :   assert (rdbk == 32'h194353) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3700   :   assert (rdbk == 32'h1b0d6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3701   :   assert (rdbk == 32'h15e377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3702   :   assert (rdbk == 32'h4bb597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3703   :   assert (rdbk == 32'hbb718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3704   :   assert (rdbk == 32'h297734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3705   :   assert (rdbk == 32'h5825b6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3706   :   assert (rdbk == 32'h2e71c6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3707   :   assert (rdbk == 32'h7b9dbd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3708   :   assert (rdbk == 32'hda6c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3709   :   assert (rdbk == 32'h154468) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3710   :   assert (rdbk == 32'h59a5e5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3711   :   assert (rdbk == 32'h682235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3712   :   assert (rdbk == 32'h6ce21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3713   :   assert (rdbk == 32'h24456b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3714   :   assert (rdbk == 32'h76b3dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3715   :   assert (rdbk == 32'h4b5710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3716   :   assert (rdbk == 32'h119d8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3717   :   assert (rdbk == 32'h75fa0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3718   :   assert (rdbk == 32'h273143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3719   :   assert (rdbk == 32'h5a2789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3720   :   assert (rdbk == 32'h4a9a98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3721   :   assert (rdbk == 32'h4ef902) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3722   :   assert (rdbk == 32'h46fb0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3723   :   assert (rdbk == 32'h189c0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3724   :   assert (rdbk == 32'h5bc20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3725   :   assert (rdbk == 32'h1bcc4f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3726   :   assert (rdbk == 32'h165399) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3727   :   assert (rdbk == 32'h625bd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3728   :   assert (rdbk == 32'h393407) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3729   :   assert (rdbk == 32'h12bc81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3730   :   assert (rdbk == 32'h33a541) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3731   :   assert (rdbk == 32'h2404e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3732   :   assert (rdbk == 32'h2d9a65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3733   :   assert (rdbk == 32'h52897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3734   :   assert (rdbk == 32'h42c763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3735   :   assert (rdbk == 32'h147670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3736   :   assert (rdbk == 32'h5ac889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3737   :   assert (rdbk == 32'h4497ff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3738   :   assert (rdbk == 32'h2ac113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3739   :   assert (rdbk == 32'h2be02e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3740   :   assert (rdbk == 32'h4d31ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3741   :   assert (rdbk == 32'h4b3417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3742   :   assert (rdbk == 32'h51182c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3743   :   assert (rdbk == 32'h253d89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3744   :   assert (rdbk == 32'h298e04) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3745   :   assert (rdbk == 32'h1550b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3746   :   assert (rdbk == 32'hce091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3747   :   assert (rdbk == 32'h7ebe85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3748   :   assert (rdbk == 32'h730c2c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3749   :   assert (rdbk == 32'h511ff2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3750   :   assert (rdbk == 32'h224dcd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3751   :   assert (rdbk == 32'h17924f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3752   :   assert (rdbk == 32'h1eea0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3753   :   assert (rdbk == 32'h17e083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3754   :   assert (rdbk == 32'h57a621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3755   :   assert (rdbk == 32'h79e657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3756   :   assert (rdbk == 32'h1e0db) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3757   :   assert (rdbk == 32'h546f1a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3758   :   assert (rdbk == 32'h9b070) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3759   :   assert (rdbk == 32'h5d862b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3760   :   assert (rdbk == 32'h62a572) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3761   :   assert (rdbk == 32'h5862d3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3762   :   assert (rdbk == 32'h326593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3763   :   assert (rdbk == 32'h44d608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3764   :   assert (rdbk == 32'h1797c6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3765   :   assert (rdbk == 32'h355faa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3766   :   assert (rdbk == 32'h3fc330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3767   :   assert (rdbk == 32'h18718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3768   :   assert (rdbk == 32'h16a2b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3769   :   assert (rdbk == 32'h1a0100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3770   :   assert (rdbk == 32'h329f1d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3771   :   assert (rdbk == 32'h256a9e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3772   :   assert (rdbk == 32'h7328ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3773   :   assert (rdbk == 32'h58d375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3774   :   assert (rdbk == 32'h580713) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3775   :   assert (rdbk == 32'h7027f0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3776   :   assert (rdbk == 32'hc561b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3777   :   assert (rdbk == 32'h594ba5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3778   :   assert (rdbk == 32'h288069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3779   :   assert (rdbk == 32'h6f179c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3780   :   assert (rdbk == 32'h291df0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3781   :   assert (rdbk == 32'h56e053) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3782   :   assert (rdbk == 32'h598995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3783   :   assert (rdbk == 32'h63b1ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3784   :   assert (rdbk == 32'h6289d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3785   :   assert (rdbk == 32'h516c9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3786   :   assert (rdbk == 32'h1c3ae2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3787   :   assert (rdbk == 32'h6e6c1e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3788   :   assert (rdbk == 32'h5111a6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3789   :   assert (rdbk == 32'h786d01) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3790   :   assert (rdbk == 32'h3ee562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3791   :   assert (rdbk == 32'h3d3aaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3792   :   assert (rdbk == 32'h1468df) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3793   :   assert (rdbk == 32'h7c2488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3794   :   assert (rdbk == 32'hc94dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3795   :   assert (rdbk == 32'h305d4f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3796   :   assert (rdbk == 32'h6b3687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3797   :   assert (rdbk == 32'h2709fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3798   :   assert (rdbk == 32'h28ef11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3799   :   assert (rdbk == 32'h3dfd5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3800   :   assert (rdbk == 32'h6996bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3801   :   assert (rdbk == 32'h5c50e6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3802   :   assert (rdbk == 32'h61acc9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3803   :   assert (rdbk == 32'hf6f9c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3804   :   assert (rdbk == 32'h5e719f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3805   :   assert (rdbk == 32'h595521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3806   :   assert (rdbk == 32'h75fd0c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3807   :   assert (rdbk == 32'h4a7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3808   :   assert (rdbk == 32'h76ec21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3809   :   assert (rdbk == 32'h39570f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3810   :   assert (rdbk == 32'h5a8c9d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3811   :   assert (rdbk == 32'h79bbaa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3812   :   assert (rdbk == 32'h4a570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3813   :   assert (rdbk == 32'h4b9b50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3814   :   assert (rdbk == 32'h738f2d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3815   :   assert (rdbk == 32'h23d51c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3816   :   assert (rdbk == 32'h74df52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3817   :   assert (rdbk == 32'h38f682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3818   :   assert (rdbk == 32'h1afa62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3819   :   assert (rdbk == 32'h73cc10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3820   :   assert (rdbk == 32'h4c1358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3821   :   assert (rdbk == 32'hb39fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3822   :   assert (rdbk == 32'h1c0835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3823   :   assert (rdbk == 32'haa37c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3824   :   assert (rdbk == 32'h244799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3825   :   assert (rdbk == 32'ha6fa8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3826   :   assert (rdbk == 32'h3caf54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3827   :   assert (rdbk == 32'hae6be) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3828   :   assert (rdbk == 32'h51639c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3829   :   assert (rdbk == 32'h18f8a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3830   :   assert (rdbk == 32'h2aedac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3831   :   assert (rdbk == 32'h3c2aac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3832   :   assert (rdbk == 32'h2f4e8d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3833   :   assert (rdbk == 32'h50198c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3834   :   assert (rdbk == 32'h41219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3835   :   assert (rdbk == 32'h42d65d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3836   :   assert (rdbk == 32'h728e08) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3837   :   assert (rdbk == 32'h29a8d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3838   :   assert (rdbk == 32'h4b5cdf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3839   :   assert (rdbk == 32'h754ce2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	// Nonce: 32'h303
	3840   :   assert (rdbk == 32'h79b387) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3841   :   assert (rdbk == 32'h6fe1dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3842   :   assert (rdbk == 32'h3219cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3843   :   assert (rdbk == 32'h5caa23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3844   :   assert (rdbk == 32'h6631b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3845   :   assert (rdbk == 32'h19d591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3846   :   assert (rdbk == 32'h416ab0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3847   :   assert (rdbk == 32'h5f6fb0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3848   :   assert (rdbk == 32'h22d66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3849   :   assert (rdbk == 32'h6a731b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3850   :   assert (rdbk == 32'h6de25a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3851   :   assert (rdbk == 32'h7534b0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3852   :   assert (rdbk == 32'h578319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3853   :   assert (rdbk == 32'h5d7805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3854   :   assert (rdbk == 32'h231264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3855   :   assert (rdbk == 32'h3447fb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3856   :   assert (rdbk == 32'h3d0b5a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3857   :   assert (rdbk == 32'h2738e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3858   :   assert (rdbk == 32'h124083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3859   :   assert (rdbk == 32'h507082) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3860   :   assert (rdbk == 32'h24f418) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3861   :   assert (rdbk == 32'h1155c9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3862   :   assert (rdbk == 32'h225499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3863   :   assert (rdbk == 32'h102101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3864   :   assert (rdbk == 32'h1507ca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3865   :   assert (rdbk == 32'h1f2ff6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3866   :   assert (rdbk == 32'h50877f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3867   :   assert (rdbk == 32'h4961e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3868   :   assert (rdbk == 32'h5a58f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3869   :   assert (rdbk == 32'h5b1479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3870   :   assert (rdbk == 32'h203a55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3871   :   assert (rdbk == 32'h232759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3872   :   assert (rdbk == 32'h1c325a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3873   :   assert (rdbk == 32'h285e5b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3874   :   assert (rdbk == 32'h150f7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3875   :   assert (rdbk == 32'h65a10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3876   :   assert (rdbk == 32'h74138c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3877   :   assert (rdbk == 32'h6be58c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3878   :   assert (rdbk == 32'h6cd6ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3879   :   assert (rdbk == 32'h3b2c7f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3880   :   assert (rdbk == 32'h5d698d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3881   :   assert (rdbk == 32'h4e3ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3882   :   assert (rdbk == 32'h5bafd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3883   :   assert (rdbk == 32'h3dda85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3884   :   assert (rdbk == 32'h2b0f0b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3885   :   assert (rdbk == 32'h33f9e8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3886   :   assert (rdbk == 32'h4f78b8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3887   :   assert (rdbk == 32'h599114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3888   :   assert (rdbk == 32'h2e0e8e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3889   :   assert (rdbk == 32'h1c5a64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3890   :   assert (rdbk == 32'h6e8f22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3891   :   assert (rdbk == 32'h22169f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3892   :   assert (rdbk == 32'h11b1ab) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3893   :   assert (rdbk == 32'h40b58a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3894   :   assert (rdbk == 32'h68f080) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3895   :   assert (rdbk == 32'hcd81e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3896   :   assert (rdbk == 32'h31933a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3897   :   assert (rdbk == 32'h6ad6d4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3898   :   assert (rdbk == 32'h32aae6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3899   :   assert (rdbk == 32'h29599b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3900   :   assert (rdbk == 32'h49d636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3901   :   assert (rdbk == 32'h5e254e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3902   :   assert (rdbk == 32'h45f7aa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3903   :   assert (rdbk == 32'h47e1d7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3904   :   assert (rdbk == 32'h3fd190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3905   :   assert (rdbk == 32'h5fb938) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3906   :   assert (rdbk == 32'h194249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3907   :   assert (rdbk == 32'h426779) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3908   :   assert (rdbk == 32'h5582c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3909   :   assert (rdbk == 32'h3ab9d5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3910   :   assert (rdbk == 32'h18089b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3911   :   assert (rdbk == 32'h535353) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3912   :   assert (rdbk == 32'h5d1022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3913   :   assert (rdbk == 32'h4c90f1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3914   :   assert (rdbk == 32'h79bebb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3915   :   assert (rdbk == 32'h78c155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3916   :   assert (rdbk == 32'h2a13f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3917   :   assert (rdbk == 32'h188d23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3918   :   assert (rdbk == 32'h4144e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3919   :   assert (rdbk == 32'h421884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3920   :   assert (rdbk == 32'h72ee7d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3921   :   assert (rdbk == 32'h5e5684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3922   :   assert (rdbk == 32'hb0a6f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3923   :   assert (rdbk == 32'h6b81d9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3924   :   assert (rdbk == 32'h3a811a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3925   :   assert (rdbk == 32'h1bad1b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3926   :   assert (rdbk == 32'h362831) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3927   :   assert (rdbk == 32'h211832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3928   :   assert (rdbk == 32'h72bc91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3929   :   assert (rdbk == 32'h5b81dc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3930   :   assert (rdbk == 32'h7e85a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3931   :   assert (rdbk == 32'h6c11fa) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3932   :   assert (rdbk == 32'h58fd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3933   :   assert (rdbk == 32'h10ce50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3934   :   assert (rdbk == 32'h7b1020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3935   :   assert (rdbk == 32'h6df0c7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3936   :   assert (rdbk == 32'h7103b9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3937   :   assert (rdbk == 32'h245f98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3938   :   assert (rdbk == 32'ha816a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3939   :   assert (rdbk == 32'h2b46ec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3940   :   assert (rdbk == 32'h73b440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3941   :   assert (rdbk == 32'h3d2f56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3942   :   assert (rdbk == 32'h5d98e6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3943   :   assert (rdbk == 32'h5658ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3944   :   assert (rdbk == 32'h477ab1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3945   :   assert (rdbk == 32'h736fb5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3946   :   assert (rdbk == 32'h5adc6e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3947   :   assert (rdbk == 32'h496b59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3948   :   assert (rdbk == 32'h188463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3949   :   assert (rdbk == 32'h30a44c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3950   :   assert (rdbk == 32'h4cbff8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3951   :   assert (rdbk == 32'h4f92cc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3952   :   assert (rdbk == 32'h7abf75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3953   :   assert (rdbk == 32'h638cfd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3954   :   assert (rdbk == 32'h724eff) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3955   :   assert (rdbk == 32'h3d88b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3956   :   assert (rdbk == 32'h2ef8d2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3957   :   assert (rdbk == 32'h309ac2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3958   :   assert (rdbk == 32'hfa9ac) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3959   :   assert (rdbk == 32'h653f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3960   :   assert (rdbk == 32'h6f1d84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3961   :   assert (rdbk == 32'h4a0a88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3962   :   assert (rdbk == 32'h4d2b06) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3963   :   assert (rdbk == 32'h83c46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3964   :   assert (rdbk == 32'h419205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3965   :   assert (rdbk == 32'h6a415b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3966   :   assert (rdbk == 32'h794c68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3967   :   assert (rdbk == 32'h44c01a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3968   :   assert (rdbk == 32'h4113dd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3969   :   assert (rdbk == 32'h486c5f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3970   :   assert (rdbk == 32'h79a7a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3971   :   assert (rdbk == 32'h7857) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3972   :   assert (rdbk == 32'h77b01f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3973   :   assert (rdbk == 32'he2ba4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3974   :   assert (rdbk == 32'h35c842) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3975   :   assert (rdbk == 32'h388815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3976   :   assert (rdbk == 32'h3d547e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3977   :   assert (rdbk == 32'h6a565a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3978   :   assert (rdbk == 32'h6e1e54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3979   :   assert (rdbk == 32'h189f11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3980   :   assert (rdbk == 32'h3aac91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3981   :   assert (rdbk == 32'h798fb2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3982   :   assert (rdbk == 32'hf854e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3983   :   assert (rdbk == 32'h13cb0f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3984   :   assert (rdbk == 32'h576295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3985   :   assert (rdbk == 32'h362ff8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3986   :   assert (rdbk == 32'h662091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3987   :   assert (rdbk == 32'h69e77f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3988   :   assert (rdbk == 32'h2f4e1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3989   :   assert (rdbk == 32'h4c5a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3990   :   assert (rdbk == 32'h14b12d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3991   :   assert (rdbk == 32'hd040a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3992   :   assert (rdbk == 32'h43ed26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3993   :   assert (rdbk == 32'h1335f6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3994   :   assert (rdbk == 32'hc6769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3995   :   assert (rdbk == 32'h4fd888) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3996   :   assert (rdbk == 32'h45b917) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3997   :   assert (rdbk == 32'h49bb57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3998   :   assert (rdbk == 32'he3b8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	3999   :   assert (rdbk == 32'h2c9cf2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4000   :   assert (rdbk == 32'h5d1e83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4001   :   assert (rdbk == 32'h26c70e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4002   :   assert (rdbk == 32'h5c6f9b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4003   :   assert (rdbk == 32'h4ab15e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4004   :   assert (rdbk == 32'h25a66d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4005   :   assert (rdbk == 32'h67b0b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4006   :   assert (rdbk == 32'h468e12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4007   :   assert (rdbk == 32'h2e313c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4008   :   assert (rdbk == 32'h4b2db0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4009   :   assert (rdbk == 32'h43906) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4010   :   assert (rdbk == 32'h126a82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4011   :   assert (rdbk == 32'h556272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4012   :   assert (rdbk == 32'h5630f3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4013   :   assert (rdbk == 32'h29ab1c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4014   :   assert (rdbk == 32'hc4425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4015   :   assert (rdbk == 32'h243da4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4016   :   assert (rdbk == 32'h7e161f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4017   :   assert (rdbk == 32'h6643c5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4018   :   assert (rdbk == 32'h10af10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4019   :   assert (rdbk == 32'h1f5f70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4020   :   assert (rdbk == 32'h4000f8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4021   :   assert (rdbk == 32'h52db10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4022   :   assert (rdbk == 32'h779946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4023   :   assert (rdbk == 32'h3693c0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4024   :   assert (rdbk == 32'h7dea36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4025   :   assert (rdbk == 32'h280e73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4026   :   assert (rdbk == 32'h3a53e3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4027   :   assert (rdbk == 32'h5e8882) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4028   :   assert (rdbk == 32'h6af0e7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4029   :   assert (rdbk == 32'h1dd75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4030   :   assert (rdbk == 32'haebb6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4031   :   assert (rdbk == 32'h7d1f05) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4032   :   assert (rdbk == 32'h783a66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4033   :   assert (rdbk == 32'h722cf5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4034   :   assert (rdbk == 32'h1a44ec) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4035   :   assert (rdbk == 32'h20d4a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4036   :   assert (rdbk == 32'h1f7c71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4037   :   assert (rdbk == 32'h253c71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4038   :   assert (rdbk == 32'h1d3084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4039   :   assert (rdbk == 32'h399d61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4040   :   assert (rdbk == 32'h6ef04f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4041   :   assert (rdbk == 32'h69496f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4042   :   assert (rdbk == 32'h5a3bda) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4043   :   assert (rdbk == 32'h5e3afb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4044   :   assert (rdbk == 32'h6998c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4045   :   assert (rdbk == 32'h45d293) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4046   :   assert (rdbk == 32'h292851) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4047   :   assert (rdbk == 32'h5c519) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4048   :   assert (rdbk == 32'h1012ae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4049   :   assert (rdbk == 32'h578ce9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4050   :   assert (rdbk == 32'h5c1ac1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4051   :   assert (rdbk == 32'h34d742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4052   :   assert (rdbk == 32'h20beca) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4053   :   assert (rdbk == 32'h56a000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4054   :   assert (rdbk == 32'h67cfe3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4055   :   assert (rdbk == 32'h2677ea) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4056   :   assert (rdbk == 32'h51ad80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4057   :   assert (rdbk == 32'h7bf217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4058   :   assert (rdbk == 32'h54a829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4059   :   assert (rdbk == 32'h359194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4060   :   assert (rdbk == 32'h321f45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4061   :   assert (rdbk == 32'h5a0f56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4062   :   assert (rdbk == 32'h1b5acc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4063   :   assert (rdbk == 32'h2f45f7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4064   :   assert (rdbk == 32'h354312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4065   :   assert (rdbk == 32'h7b875c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4066   :   assert (rdbk == 32'h5d4ae3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4067   :   assert (rdbk == 32'h416c77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4068   :   assert (rdbk == 32'h237523) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4069   :   assert (rdbk == 32'h2b453f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4070   :   assert (rdbk == 32'h1436bc) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4071   :   assert (rdbk == 32'h10a1a3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4072   :   assert (rdbk == 32'h3574bf) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4073   :   assert (rdbk == 32'h31569f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4074   :   assert (rdbk == 32'h1fab4a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4075   :   assert (rdbk == 32'h674551) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4076   :   assert (rdbk == 32'h3cbee7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4077   :   assert (rdbk == 32'h430b0d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4078   :   assert (rdbk == 32'h1f2f8f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4079   :   assert (rdbk == 32'h39e967) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4080   :   assert (rdbk == 32'h66fee4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4081   :   assert (rdbk == 32'h462499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4082   :   assert (rdbk == 32'h6e0b10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4083   :   assert (rdbk == 32'h4082a8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4084   :   assert (rdbk == 32'h10d23d) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4085   :   assert (rdbk == 32'h52a4b7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4086   :   assert (rdbk == 32'h17da74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4087   :   assert (rdbk == 32'h3e0040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4088   :   assert (rdbk == 32'h5170ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4089   :   assert (rdbk == 32'h68ad2e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4090   :   assert (rdbk == 32'h408295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4091   :   assert (rdbk == 32'h66a548) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4092   :   assert (rdbk == 32'h74c3ae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4093   :   assert (rdbk == 32'h2cd72b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4094   :   assert (rdbk == 32'h67ac0f) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	4095   :   assert (rdbk == 32'h25c181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
	
      endcase
    end

